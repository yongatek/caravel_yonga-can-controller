* NGSPICE file created from user_proj_example.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_4 abstract view
.subckt sky130_fd_sc_hd__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

.subckt user_proj_example io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ irq[0] irq[1] irq[2] la_data_in[0] la_data_in[100] la_data_in[101] la_data_in[102]
+ la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106] la_data_in[107]
+ la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112]
+ la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116] la_data_in[117]
+ la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122]
+ la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126] la_data_in[127]
+ la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17]
+ la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22]
+ la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28]
+ la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32] la_data_in[33]
+ la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38] la_data_in[39]
+ la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43] la_data_in[44]
+ la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49] la_data_in[4]
+ la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55]
+ la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5] la_data_in[60]
+ la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65] la_data_in[66]
+ la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70] la_data_in[71]
+ la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76] la_data_in[77]
+ la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81] la_data_in[82]
+ la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87] la_data_in[88]
+ la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92] la_data_in[93]
+ la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98] la_data_in[99]
+ la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] vccd1 vssd1 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3155_ _4251_/A vssd1 vssd1 vccd1 vccd1 _5544_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3086_ _3274_/B _3274_/C _3076_/Y _3079_/X _3085_/X vssd1 vssd1 vccd1 vccd1 _3086_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_39_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3988_ _3994_/A _3988_/B vssd1 vssd1 vccd1 vccd1 _3989_/A sky130_fd_sc_hd__and2_1
XANTENNA__4670__A _4824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5727_ _5736_/CLK _5727_/D vssd1 vssd1 vccd1 vccd1 _5727_/Q sky130_fd_sc_hd__dfxtp_1
X_2939_ _3321_/A _3322_/A _2944_/B _3465_/B vssd1 vssd1 vccd1 vccd1 _3053_/A sky130_fd_sc_hd__nor4b_1
XFILLER_50_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3600__C1 _3585_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5658_ _6108_/CLK _5658_/D vssd1 vssd1 vccd1 vccd1 _5658_/Q sky130_fd_sc_hd__dfxtp_1
X_5589_ _5386_/X _5580_/X _5588_/X _5586_/X vssd1 vssd1 vccd1 vccd1 _6099_/D sky130_fd_sc_hd__o211a_1
X_4609_ _5877_/Q _4579_/X _4603_/X _4608_/X vssd1 vssd1 vccd1 vccd1 _5877_/D sky130_fd_sc_hd__a22o_1
XFILLER_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4056__S _4063_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3895__S _4041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3924__A _4436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3122__A1 _4554_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output56_A _5883_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_60_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6101_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_64_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_375 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4960_ _5921_/Q _5920_/Q _5919_/Q _5918_/Q vssd1 vssd1 vccd1 vccd1 _4968_/C sky130_fd_sc_hd__and4_1
XFILLER_17_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3911_ _5233_/A _5233_/B _5236_/B vssd1 vssd1 vccd1 vccd1 _3921_/C sky130_fd_sc_hd__nor3_1
XANTENNA_clkbuf_leaf_48_wb_clk_i_A clkbuf_3_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4891_ _5951_/Q _4890_/X _4915_/S vssd1 vssd1 vccd1 vccd1 _4891_/X sky130_fd_sc_hd__mux2_1
X_3842_ _3842_/A _3842_/B vssd1 vssd1 vccd1 vccd1 _4556_/B sky130_fd_sc_hd__nand2_1
XANTENNA__5586__A _5597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3773_ _3773_/A vssd1 vssd1 vccd1 vccd1 _5706_/D sky130_fd_sc_hd__clkbuf_1
X_5512_ _5373_/X _5493_/A _5511_/X _5503_/X vssd1 vssd1 vccd1 vccd1 _6072_/D sky130_fd_sc_hd__o211a_1
XFILLER_8_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5443_ _6047_/Q _5445_/B vssd1 vssd1 vccd1 vccd1 _5443_/X sky130_fd_sc_hd__or2_1
X_5374_ _6024_/Q _5374_/B vssd1 vssd1 vccd1 vccd1 _5374_/X sky130_fd_sc_hd__or2_1
X_4325_ _3820_/A _4323_/X _5260_/A vssd1 vssd1 vccd1 vccd1 _4325_/X sky130_fd_sc_hd__o21ba_1
XFILLER_86_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4256_ _3428_/A _4252_/Y _4255_/Y _3466_/C vssd1 vssd1 vccd1 vccd1 _4256_/X sky130_fd_sc_hd__o211a_1
X_3207_ _3202_/Y _3203_/X _3204_/Y _3205_/X _3206_/Y vssd1 vssd1 vccd1 vccd1 _3214_/B
+ sky130_fd_sc_hd__o221a_1
X_4187_ _4187_/A vssd1 vssd1 vccd1 vccd1 _4200_/S sky130_fd_sc_hd__buf_2
XANTENNA__4665__A _4717_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3138_ _5738_/Q vssd1 vssd1 vccd1 vccd1 _4529_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_67_372 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3069_ _3081_/B vssd1 vssd1 vccd1 vccd1 _3266_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_27_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5496__A _6065_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3744__A _3750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4575__A _4575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5565__C1 _5556_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3654__A _3738_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3879__C1 _3432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4110_ _6113_/Q _3897_/B _4110_/S vssd1 vssd1 vccd1 vccd1 _4110_/X sky130_fd_sc_hd__mux2_1
X_5090_ _5059_/X _5080_/X _5089_/X _5087_/X vssd1 vssd1 vccd1 vccd1 _5957_/D sky130_fd_sc_hd__o211a_1
XFILLER_68_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4041_ _6098_/Q _5755_/Q _4041_/S vssd1 vssd1 vccd1 vccd1 _4041_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5992_ _5999_/CLK _5992_/D vssd1 vssd1 vccd1 vccd1 _5992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_4_wb_clk_i_A clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4943_ _5980_/Q _4928_/B _4942_/X _4940_/X vssd1 vssd1 vccd1 vccd1 _5916_/D sky130_fd_sc_hd__o211a_1
XFILLER_17_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4874_ _5965_/Q _4885_/B vssd1 vssd1 vccd1 vccd1 _4874_/X sky130_fd_sc_hd__or2_1
X_3825_ _3834_/A vssd1 vssd1 vccd1 vccd1 _3901_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3756_ _5396_/A _5702_/Q _3762_/S vssd1 vssd1 vccd1 vccd1 _3757_/B sky130_fd_sc_hd__mux2_1
XANTENNA__5308__C1 _5169_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3687_ _3770_/A vssd1 vssd1 vccd1 vccd1 _3701_/A sky130_fd_sc_hd__clkbuf_1
X_5426_ _5471_/B _5622_/B vssd1 vssd1 vccd1 vccd1 _5427_/A sky130_fd_sc_hd__or2_1
XANTENNA__3283__B _3283_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4531__B1 _4436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5357_ input7/X vssd1 vssd1 vccd1 vccd1 _5357_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_87_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5288_ _5323_/A _5301_/A _5301_/C _5288_/D vssd1 vssd1 vccd1 vccd1 _5289_/B sky130_fd_sc_hd__nand4_1
X_4308_ _5810_/Q _5809_/Q vssd1 vssd1 vccd1 vccd1 _4309_/B sky130_fd_sc_hd__nand2_1
XFILLER_87_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4239_ _4239_/A _4239_/B vssd1 vssd1 vccd1 vccd1 _4294_/A sky130_fd_sc_hd__or2_1
XFILLER_87_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3270__B1 _3269_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_proj_example_217 vssd1 vssd1 vccd1 vccd1 user_proj_example_217/HI la_data_out[124]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_206 vssd1 vssd1 vccd1 vccd1 user_proj_example_206/HI la_data_out[113]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_228 vssd1 vssd1 vccd1 vccd1 user_proj_example_228/HI wbs_dat_o[7]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_239 vssd1 vssd1 vccd1 vccd1 user_proj_example_239/HI wbs_dat_o[18]
+ sky130_fd_sc_hd__conb_1
XFILLER_2_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4590_ _6113_/Q _4588_/X _4779_/A vssd1 vssd1 vccd1 vccd1 _4590_/X sky130_fd_sc_hd__mux2_1
X_3610_ _3607_/X _3592_/X _3608_/X _3609_/X vssd1 vssd1 vccd1 vccd1 _5662_/D sky130_fd_sc_hd__o211a_1
X_3541_ _5988_/Q _4529_/A vssd1 vssd1 vccd1 vccd1 _3542_/A sky130_fd_sc_hd__nand2_1
XANTENNA__4761__A0 _6104_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3472_ _3472_/A _3017_/B vssd1 vssd1 vccd1 vccd1 _3472_/X sky130_fd_sc_hd__or2b_1
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5211_ _5220_/A _5211_/B vssd1 vssd1 vccd1 vccd1 _5212_/A sky130_fd_sc_hd__and2_1
X_5142_ _5069_/X _5125_/A _5140_/X _5141_/X vssd1 vssd1 vccd1 vccd1 _5976_/D sky130_fd_sc_hd__o211a_1
XFILLER_69_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3831__B _6121_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4816__A1 _6037_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5073_ _5953_/Q _5076_/B vssd1 vssd1 vccd1 vccd1 _5073_/X sky130_fd_sc_hd__or2_1
X_4024_ _6092_/Q _4014_/X _5750_/Q _4017_/X vssd1 vssd1 vccd1 vccd1 _4024_/X sky130_fd_sc_hd__a22o_1
XFILLER_25_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5975_ _5975_/CLK _5975_/D vssd1 vssd1 vccd1 vccd1 _5975_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4154__S _4167_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4926_ _6035_/Q _4924_/X _4925_/X _4460_/X vssd1 vssd1 vccd1 vccd1 _5909_/D sky130_fd_sc_hd__o211a_1
X_4857_ _5901_/Q _4807_/X _4853_/X _4856_/X vssd1 vssd1 vccd1 vccd1 _5901_/D sky130_fd_sc_hd__a22o_1
X_3808_ _4217_/B vssd1 vssd1 vccd1 vccd1 _3849_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4788_ _5707_/Q _5684_/Q _4797_/S vssd1 vssd1 vccd1 vccd1 _4788_/X sky130_fd_sc_hd__mux2_1
X_3739_ _3762_/S vssd1 vssd1 vccd1 vccd1 _3753_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_4_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5409_ _5461_/A vssd1 vssd1 vccd1 vccd1 _5409_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3469__A _3469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5232__A1 _5657_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3379__A _3379_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2972_ _3256_/A _3282_/B _2972_/C vssd1 vssd1 vccd1 vccd1 _2972_/X sky130_fd_sc_hd__and3_1
X_5760_ _5777_/CLK _5760_/D vssd1 vssd1 vccd1 vccd1 _5760_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5691_ _6067_/CLK _5691_/D vssd1 vssd1 vccd1 vccd1 _5691_/Q sky130_fd_sc_hd__dfxtp_1
X_4711_ _6075_/Q _4732_/B vssd1 vssd1 vccd1 vccd1 _4711_/X sky130_fd_sc_hd__or2_1
XANTENNA__5594__A _6102_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4642_ _6044_/Q _4584_/X _4610_/X _4641_/X vssd1 vssd1 vccd1 vccd1 _4642_/X sky130_fd_sc_hd__a211o_1
X_4573_ _4573_/A vssd1 vssd1 vccd1 vccd1 _5875_/D sky130_fd_sc_hd__clkbuf_1
X_3524_ _3509_/A _2955_/C _3514_/X _3523_/X vssd1 vssd1 vccd1 vccd1 _6126_/D sky130_fd_sc_hd__a31o_1
X_3455_ _3391_/A _3454_/X _3466_/D _3117_/Y _3429_/X vssd1 vssd1 vccd1 vccd1 _3455_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3842__A _3842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3386_ _3386_/A _3386_/B vssd1 vssd1 vccd1 vccd1 _3387_/A sky130_fd_sc_hd__or2_1
XFILLER_69_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5125_ _5125_/A vssd1 vssd1 vccd1 vccd1 _5125_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4149__S _4162_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5056_ _5056_/A vssd1 vssd1 vccd1 vccd1 _5056_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4007_ _4524_/A _4007_/B vssd1 vssd1 vccd1 vccd1 _4008_/A sky130_fd_sc_hd__and2_1
XFILLER_72_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5462__A1 _5393_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5958_ _5959_/CLK _5958_/D vssd1 vssd1 vccd1 vccd1 _5958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4909_ _5969_/Q _4917_/B vssd1 vssd1 vccd1 vccd1 _4909_/X sky130_fd_sc_hd__or2_1
X_5889_ _6031_/CLK _5889_/D vssd1 vssd1 vccd1 vccd1 _5889_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4612__S _4645_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4059__S _4063_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input18_A la_data_in[44] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5453__A1 _5376_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4583__A _4859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4341__A_N _5278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_3_7__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_3_7__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_16_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_14_wb_clk_i clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6122_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_3_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3240_ _5927_/Q vssd1 vssd1 vccd1 vccd1 _4986_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3171_ _3171_/A vssd1 vssd1 vccd1 vccd1 _6129_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4247__A2 _4228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5812_ _5942_/CLK _5812_/D vssd1 vssd1 vccd1 vccd1 _5812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5743_ _6131_/CLK _5743_/D vssd1 vssd1 vccd1 vccd1 _5743_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2955_ _3296_/B _5327_/B _2955_/C vssd1 vssd1 vccd1 vccd1 _2955_/X sky130_fd_sc_hd__and3_1
X_2886_ _6005_/Q vssd1 vssd1 vccd1 vccd1 _3839_/B sky130_fd_sc_hd__clkbuf_2
X_5674_ _6080_/CLK _5674_/D vssd1 vssd1 vccd1 vccd1 _5674_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4625_ _5878_/Q _4579_/X _4622_/X _4624_/Y vssd1 vssd1 vccd1 vccd1 _5878_/D sky130_fd_sc_hd__a22o_1
X_4556_ _4556_/A _4556_/B _4556_/C vssd1 vssd1 vccd1 vccd1 _4557_/S sky130_fd_sc_hd__and3_1
XANTENNA__4183__A1 _3454_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3507_ _3507_/A vssd1 vssd1 vccd1 vccd1 _3509_/B sky130_fd_sc_hd__clkinv_2
X_4487_ _4487_/A _4487_/B _4487_/C vssd1 vssd1 vccd1 vccd1 _4488_/A sky130_fd_sc_hd__or3_1
XFILLER_89_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3438_ _3438_/A _3438_/B _3833_/C vssd1 vssd1 vccd1 vccd1 _3870_/A sky130_fd_sc_hd__or3_2
X_3369_ _3380_/B _3367_/Y _3368_/X _3291_/B vssd1 vssd1 vccd1 vccd1 _3369_/X sky130_fd_sc_hd__a2bb2o_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5108_ _5045_/X _5104_/X _5107_/X _5098_/X vssd1 vssd1 vccd1 vccd1 _5963_/D sky130_fd_sc_hd__o211a_1
XFILLER_72_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6088_ _6088_/CLK _6088_/D vssd1 vssd1 vccd1 vccd1 _6088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5039_ _5944_/Q _5038_/A _5025_/B vssd1 vssd1 vccd1 vccd1 _5039_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_82_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3747__A _3750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4578__A _4858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput53 _5880_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[67] sky130_fd_sc_hd__buf_2
Xoutput64 _5891_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[78] sky130_fd_sc_hd__buf_2
Xoutput75 _5902_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[89] sky130_fd_sc_hd__buf_2
XFILLER_48_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_38_wb_clk_i_A clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4237__A_N _4327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_370 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4410_ _5839_/Q _4409_/X _4417_/S vssd1 vssd1 vccd1 vccd1 _4411_/A sky130_fd_sc_hd__mux2_1
X_5390_ _6028_/Q _5399_/B vssd1 vssd1 vccd1 vccd1 _5390_/X sky130_fd_sc_hd__or2_1
X_4341_ _5278_/A _6041_/Q vssd1 vssd1 vccd1 vccd1 _4341_/X sky130_fd_sc_hd__and2b_1
X_4272_ _4970_/A _4272_/B _4272_/C vssd1 vssd1 vccd1 vccd1 _4273_/A sky130_fd_sc_hd__and3_1
X_6011_ _6012_/CLK _6011_/D vssd1 vssd1 vccd1 vccd1 _6011_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3223_ _4946_/C vssd1 vssd1 vccd1 vccd1 _5012_/B sky130_fd_sc_hd__inv_2
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3154_ _4458_/A vssd1 vssd1 vccd1 vccd1 _4251_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_39_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3085_ _3081_/X _3082_/Y _3410_/A vssd1 vssd1 vccd1 vccd1 _3085_/X sky130_fd_sc_hd__o21a_1
XFILLER_39_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3987_ _5733_/Q _3964_/X _3953_/A _5732_/Q vssd1 vssd1 vccd1 vccd1 _3988_/B sky130_fd_sc_hd__a22o_1
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5726_ _5736_/CLK _5726_/D vssd1 vssd1 vccd1 vccd1 _5726_/Q sky130_fd_sc_hd__dfxtp_1
X_2938_ _3312_/C vssd1 vssd1 vccd1 vccd1 _3321_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__4162__S _4162_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2869_ _6005_/Q vssd1 vssd1 vccd1 vccd1 _3873_/B sky130_fd_sc_hd__inv_2
X_5657_ _6135_/CLK _5657_/D vssd1 vssd1 vccd1 vccd1 _5657_/Q sky130_fd_sc_hd__dfxtp_1
X_5588_ _6099_/Q _5592_/B vssd1 vssd1 vccd1 vccd1 _5588_/X sky130_fd_sc_hd__or2_1
X_4608_ _6017_/Q _4606_/X _4607_/X vssd1 vssd1 vccd1 vccd1 _4608_/X sky130_fd_sc_hd__o21a_1
X_4539_ _4970_/A _4539_/B vssd1 vssd1 vccd1 vccd1 _4549_/A sky130_fd_sc_hd__nand2_1
XFILLER_73_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4919__B1 _4716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_476 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4101__A _4170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5647__A1 _5382_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3940__A _3954_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output49_A _5874_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3910_ _5962_/Q _3061_/A _3909_/X vssd1 vssd1 vccd1 vccd1 _3910_/X sky130_fd_sc_hd__a21o_1
X_4890_ _6001_/Q _5993_/Q _4898_/S vssd1 vssd1 vccd1 vccd1 _4890_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3841_ _3841_/A _3841_/B _3841_/C _4220_/B vssd1 vssd1 vccd1 vccd1 _3842_/B sky130_fd_sc_hd__nor4_1
XFILLER_32_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3772_ _3784_/A _3772_/B vssd1 vssd1 vccd1 vccd1 _3773_/A sky130_fd_sc_hd__and2_1
X_5511_ _6072_/Q _5511_/B vssd1 vssd1 vccd1 vccd1 _5511_/X sky130_fd_sc_hd__or2_1
XFILLER_8_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5442_ _5366_/X _5427_/A _5441_/X _5435_/X vssd1 vssd1 vccd1 vccd1 _6046_/D sky130_fd_sc_hd__o211a_1
X_5373_ _5373_/A vssd1 vssd1 vccd1 vccd1 _5373_/X sky130_fd_sc_hd__clkbuf_2
X_4324_ _5257_/A _3406_/Y _3816_/B vssd1 vssd1 vccd1 vccd1 _5260_/A sky130_fd_sc_hd__a21bo_1
XFILLER_86_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4255_ _4255_/A _4255_/B vssd1 vssd1 vccd1 vccd1 _4255_/Y sky130_fd_sc_hd__nand2_1
XFILLER_67_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3206_ _6020_/Q _5939_/Q vssd1 vssd1 vccd1 vccd1 _3206_/Y sky130_fd_sc_hd__xnor2_1
X_4186_ _5948_/Q _5797_/Q _4196_/S vssd1 vssd1 vccd1 vccd1 _4186_/X sky130_fd_sc_hd__mux2_1
X_3137_ _4562_/B _3129_/X _3135_/X _3999_/A vssd1 vssd1 vccd1 vccd1 _5737_/D sky130_fd_sc_hd__a211o_1
XFILLER_67_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4157__S _4167_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3068_ _5856_/Q vssd1 vssd1 vccd1 vccd1 _3081_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_63_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3297__A _3317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5709_ _5996_/CLK _5709_/D vssd1 vssd1 vccd1 vccd1 _5709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4301__A1 _4233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3654__B _5174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3879__B1 _4466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3092__D _3272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4040_ _4040_/A vssd1 vssd1 vccd1 vccd1 _5755_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_151 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5253__C1 _4288_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5991_ _5999_/CLK _5991_/D vssd1 vssd1 vccd1 vccd1 _5991_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5597__A _5597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4942_ _5916_/Q _4942_/B vssd1 vssd1 vccd1 vccd1 _4942_/X sky130_fd_sc_hd__or2_1
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4873_ _5957_/Q _4872_/X _4873_/S vssd1 vssd1 vccd1 vccd1 _4873_/X sky130_fd_sc_hd__mux2_1
X_3824_ _3824_/A _4002_/A _3840_/B _3824_/D vssd1 vssd1 vccd1 vccd1 _3834_/A sky130_fd_sc_hd__and4_1
X_3755_ _3755_/A vssd1 vssd1 vccd1 vccd1 _5701_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3686_ _4251_/A vssd1 vssd1 vccd1 vccd1 _3770_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3564__B _3564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5425_ _3617_/X _5404_/A _5424_/X _5420_/X vssd1 vssd1 vccd1 vccd1 _6040_/D sky130_fd_sc_hd__o211a_1
X_5356_ _5353_/X _5347_/X _5354_/Y _5355_/X vssd1 vssd1 vccd1 vccd1 _6018_/D sky130_fd_sc_hd__o211a_1
X_5287_ _5287_/A _5287_/B _5287_/C _5287_/D vssd1 vssd1 vccd1 vccd1 _5287_/X sky130_fd_sc_hd__or4_1
X_4307_ _4307_/A _4307_/B vssd1 vssd1 vccd1 vccd1 _4307_/Y sky130_fd_sc_hd__nor2_1
XFILLER_59_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3098__A1 _3481_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4238_ _6129_/Q vssd1 vssd1 vccd1 vccd1 _4239_/A sky130_fd_sc_hd__inv_2
XANTENNA__3098__B2 _3159_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4295__B1 _3723_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_535 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4169_ _5661_/Q _5792_/Q _4179_/S vssd1 vssd1 vccd1 vccd1 _4169_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4615__S _5603_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_proj_example_218 vssd1 vssd1 vccd1 vccd1 user_proj_example_218/HI la_data_out[125]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_207 vssd1 vssd1 vccd1 vccd1 user_proj_example_207/HI la_data_out[114]
+ sky130_fd_sc_hd__conb_1
XFILLER_11_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xuser_proj_example_229 vssd1 vssd1 vccd1 vccd1 user_proj_example_229/HI wbs_dat_o[8]
+ sky130_fd_sc_hd__conb_1
XFILLER_78_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input48_A wbs_we_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4586__A _4870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3490__A _4113_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_39_wb_clk_i clkbuf_3_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5975_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_3_5__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3540_ _4545_/A _5868_/Q _4541_/A _4534_/A vssd1 vssd1 vccd1 vccd1 _3540_/X sky130_fd_sc_hd__or4_1
X_3471_ _5279_/A _3469_/B _3007_/X _3293_/A _3854_/A vssd1 vssd1 vccd1 vccd1 _3472_/A
+ sky130_fd_sc_hd__o32a_1
X_5210_ _5059_/A _5999_/Q _5216_/S vssd1 vssd1 vccd1 vccd1 _5211_/B sky130_fd_sc_hd__mux2_1
XFILLER_69_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5141_ _5141_/A vssd1 vssd1 vccd1 vccd1 _5141_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5072_ _5072_/A vssd1 vssd1 vccd1 vccd1 _5072_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4023_ _4023_/A vssd1 vssd1 vccd1 vccd1 _5750_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5474__C1 _5461_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5974_ _5974_/CLK _5974_/D vssd1 vssd1 vccd1 vccd1 _5974_/Q sky130_fd_sc_hd__dfxtp_1
X_4925_ _5909_/Q _4942_/B vssd1 vssd1 vccd1 vccd1 _4925_/X sky130_fd_sc_hd__or2_1
X_4856_ _5979_/Q _4854_/X _4855_/X vssd1 vssd1 vccd1 vccd1 _4856_/X sky130_fd_sc_hd__o21a_1
X_3807_ _4220_/A _3928_/A vssd1 vssd1 vccd1 vccd1 _4217_/B sky130_fd_sc_hd__nor2_1
XANTENNA__3575__A _5622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4787_ _5894_/Q _4756_/X _4785_/X _4786_/X vssd1 vssd1 vccd1 vccd1 _5894_/D sky130_fd_sc_hd__a22o_1
X_3738_ _3738_/A _5201_/A vssd1 vssd1 vccd1 vccd1 _3762_/S sky130_fd_sc_hd__nand2_1
X_3669_ _5393_/A _5678_/Q _3669_/S vssd1 vssd1 vccd1 vccd1 _3670_/B sky130_fd_sc_hd__mux2_1
X_5408_ _5408_/A vssd1 vssd1 vccd1 vccd1 _5461_/A sky130_fd_sc_hd__clkbuf_2
X_5339_ _6068_/Q _6015_/Q _5339_/S vssd1 vssd1 vccd1 vccd1 _5339_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_6__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5836_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_55_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5232__A2 _3061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4743__A1 _6054_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2971_ _3321_/A _3438_/B _3288_/C vssd1 vssd1 vccd1 vccd1 _3282_/B sky130_fd_sc_hd__and3_1
XFILLER_61_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5690_ _6067_/CLK _5690_/D vssd1 vssd1 vccd1 vccd1 _5690_/Q sky130_fd_sc_hd__dfxtp_1
X_4710_ _6099_/Q _4709_/X _4720_/S vssd1 vssd1 vccd1 vccd1 _4710_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4641_ _4611_/X _4638_/X _4640_/X _4620_/X vssd1 vssd1 vccd1 vccd1 _4641_/X sky130_fd_sc_hd__o211a_1
X_4572_ _5186_/A _4572_/B vssd1 vssd1 vccd1 vccd1 _4573_/A sky130_fd_sc_hd__and2_1
XANTENNA__3826__C _3826_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3523_ _5278_/A _3519_/X _3520_/X _3505_/C _3522_/X vssd1 vssd1 vccd1 vccd1 _3523_/X
+ sky130_fd_sc_hd__a221o_1
X_3454_ _4283_/A vssd1 vssd1 vccd1 vccd1 _3454_/X sky130_fd_sc_hd__clkbuf_4
X_3385_ _4409_/S _3369_/X _3377_/X _3384_/X vssd1 vssd1 vccd1 vccd1 _3386_/B sky130_fd_sc_hd__a211o_1
XFILLER_57_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5124_ _5469_/B _5148_/B vssd1 vssd1 vccd1 vccd1 _5125_/A sky130_fd_sc_hd__or2_1
XFILLER_29_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5055_ _5045_/X _5050_/X _5054_/X _5043_/X vssd1 vssd1 vccd1 vccd1 _5947_/D sky130_fd_sc_hd__o211a_1
X_4006_ _5746_/Q _3927_/Y _4006_/S vssd1 vssd1 vccd1 vccd1 _4007_/B sky130_fd_sc_hd__mux2_1
XFILLER_65_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5957_ _5959_/CLK _5957_/D vssd1 vssd1 vccd1 vccd1 _5957_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4908_ _5961_/Q _4907_/X _4916_/S vssd1 vssd1 vccd1 vccd1 _4908_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5888_ _6031_/CLK _5888_/D vssd1 vssd1 vccd1 vccd1 _5888_/Q sky130_fd_sc_hd__dfxtp_1
X_4839_ _5712_/Q _5689_/Q _4848_/S vssd1 vssd1 vccd1 vccd1 _4839_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4725__A1 _6028_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_438 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_28_wb_clk_i_A clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_43_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5610__C1 _5597_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3927__B _6121_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_54_wb_clk_i clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _5892_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3170_ _3632_/A _3170_/B vssd1 vssd1 vccd1 vccd1 _3171_/A sky130_fd_sc_hd__and2_1
XFILLER_86_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3455__A1 _3391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5811_ _5942_/CLK _5811_/D vssd1 vssd1 vccd1 vccd1 _5811_/Q sky130_fd_sc_hd__dfxtp_1
X_5742_ _5874_/CLK _5742_/D vssd1 vssd1 vccd1 vccd1 _5742_/Q sky130_fd_sc_hd__dfxtp_1
X_2954_ _5241_/B _3836_/A vssd1 vssd1 vccd1 vccd1 _2955_/C sky130_fd_sc_hd__nor2_2
X_2885_ _3071_/A _2885_/B vssd1 vssd1 vccd1 vccd1 _2885_/Y sky130_fd_sc_hd__nor2_1
X_5673_ _6077_/CLK _5673_/D vssd1 vssd1 vccd1 vccd1 _5673_/Q sky130_fd_sc_hd__dfxtp_1
X_4624_ _5354_/A _4602_/X _4623_/X vssd1 vssd1 vccd1 vccd1 _4624_/Y sky130_fd_sc_hd__a21oi_1
X_4555_ _5254_/A _4555_/B _4555_/C vssd1 vssd1 vccd1 vccd1 _4556_/A sky130_fd_sc_hd__nor3_1
X_3506_ _3255_/X _4409_/S _3504_/X _3505_/X vssd1 vssd1 vccd1 vccd1 _6124_/D sky130_fd_sc_hd__a31o_1
X_4486_ _5870_/Q _5869_/Q _4534_/A _4534_/B vssd1 vssd1 vccd1 vccd1 _4487_/C sky130_fd_sc_hd__or4b_1
XFILLER_89_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3437_ _3424_/X _2972_/X _3300_/A _3434_/Y _3436_/Y vssd1 vssd1 vccd1 vccd1 _3437_/X
+ sky130_fd_sc_hd__a221o_1
X_3368_ _3897_/A _3493_/A _3368_/C vssd1 vssd1 vccd1 vccd1 _3368_/X sky130_fd_sc_hd__and3_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5107_ _5963_/Q _5116_/B vssd1 vssd1 vccd1 vccd1 _5107_/X sky130_fd_sc_hd__or2_1
X_3299_ _4470_/A _4283_/B _3829_/D _3380_/B vssd1 vssd1 vccd1 vccd1 _3299_/X sky130_fd_sc_hd__or4_1
X_6087_ _6087_/CLK _6087_/D vssd1 vssd1 vccd1 vccd1 _6087_/Q sky130_fd_sc_hd__dfxtp_1
X_5038_ _5038_/A _5038_/B vssd1 vssd1 vccd1 vccd1 _5943_/D sky130_fd_sc_hd__nor2_1
XFILLER_25_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4859__A _4859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput65 _5892_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[79] sky130_fd_sc_hd__buf_2
Xoutput76 _5903_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[90] sky130_fd_sc_hd__buf_2
Xoutput54 _5881_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[68] sky130_fd_sc_hd__buf_2
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_511 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input30_A la_data_in[55] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_40 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3938__A _3938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5362__A1 _5360_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4340_ _4340_/A vssd1 vssd1 vccd1 vccd1 _5818_/D sky130_fd_sc_hd__clkbuf_1
X_4271_ _5807_/Q _4275_/C vssd1 vssd1 vccd1 vccd1 _4272_/C sky130_fd_sc_hd__xor2_1
X_6010_ _6012_/CLK _6010_/D vssd1 vssd1 vccd1 vccd1 _6010_/Q sky130_fd_sc_hd__dfxtp_1
X_3222_ _5011_/B _4942_/B _3219_/X _3221_/X vssd1 vssd1 vccd1 vccd1 _5854_/D sky130_fd_sc_hd__o31a_1
X_3153_ _3375_/B vssd1 vssd1 vccd1 vccd1 _4458_/A sky130_fd_sc_hd__clkinv_2
XFILLER_39_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3084_ _4466_/A vssd1 vssd1 vccd1 vccd1 _3410_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_50_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3986_ _3999_/A _3986_/B vssd1 vssd1 vccd1 vccd1 _5732_/D sky130_fd_sc_hd__nor2_1
XFILLER_50_455 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2937_ _3466_/C _3047_/A _5301_/B vssd1 vssd1 vccd1 vccd1 _5289_/A sky130_fd_sc_hd__o21ai_1
X_5725_ _5736_/CLK _5725_/D vssd1 vssd1 vccd1 vccd1 _5725_/Q sky130_fd_sc_hd__dfxtp_1
X_5656_ _6135_/CLK _5656_/D vssd1 vssd1 vccd1 vccd1 _5656_/Q sky130_fd_sc_hd__dfxtp_1
X_2868_ _3459_/D vssd1 vssd1 vccd1 vccd1 _3071_/A sky130_fd_sc_hd__buf_2
X_4607_ _4607_/A vssd1 vssd1 vccd1 vccd1 _4607_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5587_ _5382_/X _5580_/X _5585_/X _5586_/X vssd1 vssd1 vccd1 vccd1 _6098_/D sky130_fd_sc_hd__o211a_1
XANTENNA__3583__A _5657_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4538_ _4562_/A _4538_/B _4527_/X vssd1 vssd1 vccd1 vccd1 _4539_/B sky130_fd_sc_hd__or3b_1
XFILLER_77_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4469_ _5954_/Q _3061_/A _4468_/X vssd1 vssd1 vccd1 vccd1 _4469_/X sky130_fd_sc_hd__a21o_1
XFILLER_77_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5041__B1 _3221_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_488 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3668__A _3668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3840_ _4002_/A _3840_/B vssd1 vssd1 vccd1 vccd1 _4220_/B sky130_fd_sc_hd__nand2_1
X_3771_ _3598_/A _5706_/Q _3780_/S vssd1 vssd1 vccd1 vccd1 _3772_/B sky130_fd_sc_hd__mux2_1
X_5510_ _5369_/X _5493_/A _5509_/X _5503_/X vssd1 vssd1 vccd1 vccd1 _6071_/D sky130_fd_sc_hd__o211a_1
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5441_ _6046_/Q _5445_/B vssd1 vssd1 vccd1 vccd1 _5441_/X sky130_fd_sc_hd__or2_1
X_5372_ _5369_/X _5354_/B _5370_/X _5371_/X vssd1 vssd1 vccd1 vccd1 _6023_/D sky130_fd_sc_hd__o211a_1
X_4323_ _4294_/B _4320_/Y _4321_/X _4294_/A _4322_/Y vssd1 vssd1 vccd1 vccd1 _4323_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_59_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4254_ _3843_/B _3482_/B _4253_/X vssd1 vssd1 vccd1 vccd1 _4255_/B sky130_fd_sc_hd__a21oi_1
X_3205_ _6022_/Q _5941_/Q vssd1 vssd1 vccd1 vccd1 _3205_/X sky130_fd_sc_hd__and2_1
X_4185_ _4185_/A vssd1 vssd1 vccd1 vccd1 _5797_/D sky130_fd_sc_hd__clkbuf_1
X_3136_ _3547_/A vssd1 vssd1 vccd1 vccd1 _3999_/A sky130_fd_sc_hd__buf_4
XFILLER_67_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3067_ _3067_/A vssd1 vssd1 vccd1 vccd1 _3423_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3578__A _5622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5574__A1 _5366_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3969_ _5728_/Q _3964_/X _3945_/X _5727_/Q vssd1 vssd1 vccd1 vccd1 _3970_/B sky130_fd_sc_hd__a22o_1
X_5708_ _6085_/CLK _5708_/D vssd1 vssd1 vccd1 vccd1 _5708_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5639_ _5366_/X _5623_/A _5637_/X _5638_/X vssd1 vssd1 vccd1 vccd1 _6118_/D sky130_fd_sc_hd__o211a_1
XFILLER_77_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5565__A1 _5353_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output61_A _5888_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5990_ _5999_/CLK _5990_/D vssd1 vssd1 vccd1 vccd1 _5990_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3803__A1 _4409_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4941_ _5979_/Q _4928_/B _4939_/Y _4940_/X vssd1 vssd1 vccd1 vccd1 _5915_/D sky130_fd_sc_hd__o211a_1
XFILLER_52_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4872_ _5949_/Q _4871_/X _4872_/S vssd1 vssd1 vccd1 vccd1 _4872_/X sky130_fd_sc_hd__mux2_1
X_3823_ _2858_/A _5754_/Q _3820_/Y _3822_/X vssd1 vssd1 vccd1 vccd1 _3823_/X sky130_fd_sc_hd__o31a_1
XFILLER_20_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_9_wb_clk_i _5813_/CLK vssd1 vssd1 vccd1 vccd1 _6005_/CLK sky130_fd_sc_hd__clkbuf_16
X_3754_ _3768_/A _3754_/B vssd1 vssd1 vccd1 vccd1 _3755_/A sky130_fd_sc_hd__and2_1
XANTENNA__3845__B _4438_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3685_ _3685_/A vssd1 vssd1 vccd1 vccd1 _5682_/D sky130_fd_sc_hd__clkbuf_1
X_5424_ _6040_/Q _5424_/B vssd1 vssd1 vccd1 vccd1 _5424_/X sky130_fd_sc_hd__or2_1
XFILLER_87_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5355_ _5391_/A vssd1 vssd1 vccd1 vccd1 _5355_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5286_ _5297_/B _5297_/C vssd1 vssd1 vccd1 vccd1 _5288_/D sky130_fd_sc_hd__or2_1
X_4306_ _4306_/A _4306_/B _4306_/C _4306_/D vssd1 vssd1 vccd1 vccd1 _4307_/B sky130_fd_sc_hd__or4_1
XFILLER_59_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4237_ _4327_/A _4241_/A _4237_/C vssd1 vssd1 vccd1 vccd1 _4329_/B sky130_fd_sc_hd__and3b_1
XFILLER_55_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_5__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_3_5__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_28_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4168_ _4168_/A vssd1 vssd1 vccd1 vccd1 _5792_/D sky130_fd_sc_hd__clkbuf_1
X_3119_ _5245_/A vssd1 vssd1 vccd1 vccd1 _5243_/B sky130_fd_sc_hd__clkbuf_2
X_4099_ _5959_/Q _5772_/Q _4110_/S vssd1 vssd1 vccd1 vccd1 _4099_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3270__A2 _3891_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xuser_proj_example_208 vssd1 vssd1 vccd1 vccd1 user_proj_example_208/HI la_data_out[115]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_219 vssd1 vssd1 vccd1 vccd1 user_proj_example_219/HI la_data_out[126]
+ sky130_fd_sc_hd__conb_1
XANTENNA__4507__C1 _4460_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4286__A1 _3839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_536 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4038__A1 _6097_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3011__A _3836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2850__A _3038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3470_ _3469_/A _3434_/A _2983_/B _3469_/X vssd1 vssd1 vccd1 vccd1 _3470_/X sky130_fd_sc_hd__o31a_1
XFILLER_6_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3681__A _3765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3721__B1 _3999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5140_ _5976_/Q _5145_/B vssd1 vssd1 vccd1 vccd1 _5140_/X sky130_fd_sc_hd__or2_1
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5071_ _5069_/X _5050_/A _5070_/X _5067_/X vssd1 vssd1 vccd1 vccd1 _5952_/D sky130_fd_sc_hd__o211a_1
XFILLER_84_428 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4022_ _5750_/Q _4021_/X _4028_/S vssd1 vssd1 vccd1 vccd1 _4023_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5401__A _5401_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5973_ _5974_/CLK _5973_/D vssd1 vssd1 vccd1 vccd1 _5973_/Q sky130_fd_sc_hd__dfxtp_1
X_4924_ _4944_/B vssd1 vssd1 vccd1 vccd1 _4924_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4855_ _4855_/A vssd1 vssd1 vccd1 vccd1 _4855_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3806_ _3806_/A vssd1 vssd1 vccd1 vccd1 _5714_/D sky130_fd_sc_hd__clkbuf_1
X_4786_ _6034_/Q _4744_/X _4745_/X vssd1 vssd1 vccd1 vccd1 _4786_/X sky130_fd_sc_hd__o21a_1
XANTENNA__3575__B _5579_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3737_ _3737_/A vssd1 vssd1 vccd1 vccd1 _5696_/D sky130_fd_sc_hd__clkbuf_1
X_3668_ _3668_/A vssd1 vssd1 vccd1 vccd1 _3684_/A sky130_fd_sc_hd__clkbuf_1
X_3599_ _5659_/Q _3608_/B vssd1 vssd1 vccd1 vccd1 _3599_/X sky130_fd_sc_hd__or2_1
XANTENNA__3591__A _5622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5407_ _6033_/Q _5417_/B vssd1 vssd1 vccd1 vccd1 _5407_/X sky130_fd_sc_hd__or2_1
X_5338_ _5338_/A vssd1 vssd1 vccd1 vccd1 _6015_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2919__B _2941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5269_ _5269_/A _5269_/B _5269_/C _5287_/D vssd1 vssd1 vccd1 vccd1 _5269_/X sky130_fd_sc_hd__or4_1
XFILLER_75_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_18_wb_clk_i_A _5836_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4626__S _4645_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_57_wb_clk_i_A clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_78_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2970_ _3465_/C vssd1 vssd1 vccd1 vccd1 _3438_/B sky130_fd_sc_hd__inv_2
XFILLER_61_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4640_ _6068_/Q _4683_/B vssd1 vssd1 vccd1 vccd1 _4640_/X sky130_fd_sc_hd__or2_1
XANTENNA__3395__B _3826_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4571_ _4567_/Y _3556_/A _4575_/B _5875_/Q vssd1 vssd1 vccd1 vccd1 _4572_/B sky130_fd_sc_hd__a2bb2o_1
X_3522_ _3522_/A _3522_/B _3522_/C vssd1 vssd1 vccd1 vccd1 _3522_/X sky130_fd_sc_hd__and3_1
XFILLER_89_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3453_ _3433_/Y _3437_/X _3441_/X _3452_/X _3158_/A vssd1 vssd1 vccd1 vccd1 _3489_/A
+ sky130_fd_sc_hd__o41a_1
XFILLER_69_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3384_ _4206_/A _4450_/B _3380_/Y _4366_/A _3423_/B vssd1 vssd1 vccd1 vccd1 _3384_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_69_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5123_ _5075_/X _5104_/A _5122_/X _5114_/X vssd1 vssd1 vccd1 vccd1 _5970_/D sky130_fd_sc_hd__o211a_1
X_5054_ _5947_/Q _5066_/B vssd1 vssd1 vccd1 vccd1 _5054_/X sky130_fd_sc_hd__or2_1
X_4005_ _4450_/B _4001_/Y _4452_/S vssd1 vssd1 vccd1 vccd1 _4006_/S sky130_fd_sc_hd__a21o_1
XFILLER_65_483 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4970__A _4970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5956_ _5959_/CLK _5956_/D vssd1 vssd1 vccd1 vccd1 _5956_/Q sky130_fd_sc_hd__dfxtp_1
X_5887_ _6031_/CLK _5887_/D vssd1 vssd1 vccd1 vccd1 _5887_/Q sky130_fd_sc_hd__dfxtp_1
X_4907_ _5953_/Q _4906_/X _4915_/S vssd1 vssd1 vccd1 vccd1 _4907_/X sky130_fd_sc_hd__mux2_1
X_4838_ _5899_/Q _4807_/X _4836_/X _4837_/X vssd1 vssd1 vccd1 vccd1 _5899_/D sky130_fd_sc_hd__a22o_1
X_4769_ _5705_/Q _5682_/Q _4797_/S vssd1 vssd1 vccd1 vccd1 _4769_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4210__A _4210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4864__B _4885_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4110__A0 _6113_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_23_wb_clk_i clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5926_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_66_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3455__A2 _3454_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4652__A1 _5881_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5810_ _5942_/CLK _5810_/D vssd1 vssd1 vccd1 vccd1 _5810_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5741_ _6121_/CLK _5741_/D vssd1 vssd1 vccd1 vccd1 _5741_/Q sky130_fd_sc_hd__dfxtp_1
X_2953_ _3296_/A vssd1 vssd1 vccd1 vccd1 _5241_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_62_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2884_ _3873_/B _3304_/B vssd1 vssd1 vccd1 vccd1 _2885_/B sky130_fd_sc_hd__nand2_1
XFILLER_30_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5672_ _6027_/CLK _5672_/D vssd1 vssd1 vccd1 vccd1 _5672_/Q sky130_fd_sc_hd__dfxtp_1
X_4623_ _4858_/A vssd1 vssd1 vccd1 vccd1 _4623_/X sky130_fd_sc_hd__clkbuf_2
X_4554_ _5665_/Q _4553_/X _4554_/S vssd1 vssd1 vccd1 vccd1 _4554_/X sky130_fd_sc_hd__mux2_1
X_3505_ _3668_/A _3935_/C _3505_/C vssd1 vssd1 vccd1 vccd1 _3505_/X sky130_fd_sc_hd__and3_1
X_4485_ _5865_/Q vssd1 vssd1 vccd1 vccd1 _4534_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3436_ _3469_/B _3293_/A _4259_/B _3435_/X vssd1 vssd1 vccd1 vccd1 _3436_/Y sky130_fd_sc_hd__o31ai_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3367_ _3494_/A _3891_/B vssd1 vssd1 vccd1 vccd1 _3367_/Y sky130_fd_sc_hd__nand2_1
XFILLER_85_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6086_ _6087_/CLK _6086_/D vssd1 vssd1 vccd1 vccd1 _6086_/Q sky130_fd_sc_hd__dfxtp_1
X_5106_ _5122_/B vssd1 vssd1 vccd1 vccd1 _5116_/B sky130_fd_sc_hd__clkbuf_1
X_3298_ _3298_/A _5245_/A _3836_/A _3298_/D vssd1 vssd1 vccd1 vccd1 _3380_/B sky130_fd_sc_hd__or4_2
X_5037_ _5943_/Q _5035_/A _5020_/X vssd1 vssd1 vccd1 vccd1 _5038_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__4643__A1 _6020_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5939_ _5944_/CLK _5939_/D vssd1 vssd1 vccd1 vccd1 _5939_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3603__C1 _3585_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3466__D _3466_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput66 _5893_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[80] sky130_fd_sc_hd__buf_2
Xoutput55 _5882_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[69] sky130_fd_sc_hd__buf_2
Xoutput77 _5904_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[91] sky130_fd_sc_hd__buf_2
XFILLER_76_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input23_A la_data_in[49] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4634__A1 _6019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3954__A _3954_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4270_ _4270_/A _4270_/B _4270_/C _4228_/X vssd1 vssd1 vccd1 vccd1 _4272_/B sky130_fd_sc_hd__or4b_1
X_3221_ _5638_/A vssd1 vssd1 vccd1 vccd1 _3221_/X sky130_fd_sc_hd__clkbuf_4
X_3152_ _3139_/Y _5284_/A _3149_/X _4462_/S vssd1 vssd1 vccd1 vccd1 _5738_/D sky130_fd_sc_hd__o31ai_1
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3083_ _5241_/B vssd1 vssd1 vccd1 vccd1 _4466_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__4625__A1 _5878_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3985_ _5732_/Q _3932_/A _3984_/X vssd1 vssd1 vccd1 vccd1 _3986_/B sky130_fd_sc_hd__a21oi_1
X_2936_ _2936_/A _3317_/A vssd1 vssd1 vccd1 vccd1 _5301_/B sky130_fd_sc_hd__or2_1
X_5724_ _5736_/CLK _5724_/D vssd1 vssd1 vccd1 vccd1 _5724_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2867_ _3842_/A vssd1 vssd1 vccd1 vccd1 _3459_/D sky130_fd_sc_hd__clkbuf_2
X_5655_ _5396_/X _3576_/A _5654_/X _5172_/X vssd1 vssd1 vccd1 vccd1 _6138_/D sky130_fd_sc_hd__o211a_1
X_4606_ _5379_/B vssd1 vssd1 vccd1 vccd1 _4606_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5586_ _5597_/A vssd1 vssd1 vccd1 vccd1 _5586_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4537_ _4537_/A vssd1 vssd1 vccd1 vccd1 _5866_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4561__B1 _3245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4468_ _3917_/A _3462_/X _4467_/X _3331_/X vssd1 vssd1 vccd1 vccd1 _4468_/X sky130_fd_sc_hd__o211a_1
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3419_ _5854_/Q _3218_/X _3418_/Y vssd1 vssd1 vccd1 vccd1 _3420_/B sky130_fd_sc_hd__a21oi_1
X_4399_ _6059_/Q _3357_/X _4399_/S vssd1 vssd1 vccd1 vccd1 _4400_/A sky130_fd_sc_hd__mux2_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6138_ _6138_/CLK _6138_/D vssd1 vssd1 vccd1 vccd1 _6138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3104__A _5250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6069_ _6091_/CLK _6069_/D vssd1 vssd1 vccd1 vccd1 _6069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4919__A2 _4706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5501__C1 _5488_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3014__A _3038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2853__A _3272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3770_ _3770_/A vssd1 vssd1 vccd1 vccd1 _3784_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_12_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5440_ _5363_/X _5427_/X _5439_/X _5435_/X vssd1 vssd1 vccd1 vccd1 _6045_/D sky130_fd_sc_hd__o211a_1
XFILLER_66_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5371_ _5391_/A vssd1 vssd1 vccd1 vccd1 _5371_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4322_ _4322_/A _4322_/B vssd1 vssd1 vccd1 vccd1 _4322_/Y sky130_fd_sc_hd__nand2_1
X_4253_ _3052_/A _3826_/C _3427_/C _4438_/B vssd1 vssd1 vccd1 vccd1 _4253_/X sky130_fd_sc_hd__o211a_1
XFILLER_4_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_128 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3204_ _6022_/Q _5941_/Q vssd1 vssd1 vccd1 vccd1 _3204_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4846__A1 _6040_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4184_ _5797_/Q _4183_/X _4184_/S vssd1 vssd1 vccd1 vccd1 _4185_/A sky130_fd_sc_hd__mux2_1
X_3135_ _3135_/A _4562_/A _3135_/C vssd1 vssd1 vccd1 vccd1 _3135_/X sky130_fd_sc_hd__and3_1
XFILLER_55_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_3_4__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_3_4__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
X_3066_ _3373_/A _3066_/B vssd1 vssd1 vccd1 vccd1 _3067_/A sky130_fd_sc_hd__nand2_1
XFILLER_82_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3578__B _5581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3968_ _5188_/A vssd1 vssd1 vccd1 vccd1 _3994_/A sky130_fd_sc_hd__clkbuf_1
X_2919_ _3460_/A _2941_/A _5323_/B vssd1 vssd1 vccd1 vccd1 _3058_/A sky130_fd_sc_hd__or3_1
XFILLER_50_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5707_ _6085_/CLK _5707_/D vssd1 vssd1 vccd1 vccd1 _5707_/Q sky130_fd_sc_hd__dfxtp_1
X_3899_ _3899_/A vssd1 vssd1 vccd1 vccd1 _3899_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3594__A _5624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5638_ _5638_/A vssd1 vssd1 vccd1 vccd1 _5638_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3337__B2 _3841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5569_ _5360_/X _5559_/X _5568_/X _5556_/X vssd1 vssd1 vccd1 vccd1 _6092_/D sky130_fd_sc_hd__o211a_1
XFILLER_2_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4837__A1 _6039_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3009__A _3824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output54_A _5881_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4461__C1 _4460_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4940_ _5067_/A vssd1 vssd1 vccd1 vccd1 _4940_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4871_ _5999_/Q _5991_/Q _4898_/S vssd1 vssd1 vccd1 vccd1 _4871_/X sky130_fd_sc_hd__mux2_1
X_3822_ _3071_/A _3821_/X _6096_/Q _3331_/X vssd1 vssd1 vccd1 vccd1 _3822_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_20_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3753_ _5393_/A _5701_/Q _3753_/S vssd1 vssd1 vccd1 vccd1 _3754_/B sky130_fd_sc_hd__mux2_1
XFILLER_9_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3684_ _3684_/A _3684_/B vssd1 vssd1 vccd1 vccd1 _3685_/A sky130_fd_sc_hd__and2_1
X_5423_ _3614_/X _5404_/A _5422_/X _5420_/X vssd1 vssd1 vccd1 vccd1 _6039_/D sky130_fd_sc_hd__o211a_1
X_5354_ _5354_/A _5354_/B vssd1 vssd1 vccd1 vccd1 _5354_/Y sky130_fd_sc_hd__nand2_1
X_4305_ _3275_/X _3497_/X _4294_/B vssd1 vssd1 vccd1 vccd1 _4306_/D sky130_fd_sc_hd__a21oi_1
X_5285_ _5285_/A vssd1 vssd1 vccd1 vccd1 _5323_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5134__A _5973_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4236_ _4236_/A _5252_/B vssd1 vssd1 vccd1 vccd1 _4327_/A sky130_fd_sc_hd__or2_2
X_4167_ _5792_/Q _4166_/X _4167_/S vssd1 vssd1 vccd1 vccd1 _4168_/A sky130_fd_sc_hd__mux2_1
X_3118_ _3161_/A _3118_/B vssd1 vssd1 vccd1 vccd1 _3118_/Y sky130_fd_sc_hd__nand2_1
XFILLER_55_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4098_ _4098_/A vssd1 vssd1 vccd1 vccd1 _5772_/D sky130_fd_sc_hd__clkbuf_1
X_3049_ _3049_/A _5851_/Q vssd1 vssd1 vccd1 vccd1 _3427_/C sky130_fd_sc_hd__xnor2_1
XFILLER_55_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4184__S _4184_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_proj_example_209 vssd1 vssd1 vccd1 vccd1 user_proj_example_209/HI la_data_out[116]
+ sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_leaf_47_wb_clk_i_A clkbuf_3_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_78_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4883__A _4883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4038__A2 _3491_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3246__B1 _3245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_48_wb_clk_i clkbuf_3_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6085_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__3549__B2 _3255_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3681__B _5174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3721__A1 _4575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5070_ _5952_/Q _5076_/B vssd1 vssd1 vccd1 vccd1 _5070_/X sky130_fd_sc_hd__or2_1
XFILLER_84_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4021_ _6091_/Q _4014_/X _5749_/Q _4017_/X vssd1 vssd1 vccd1 vccd1 _4021_/X sky130_fd_sc_hd__a22o_1
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5972_ _5974_/CLK _5972_/D vssd1 vssd1 vccd1 vccd1 _5972_/Q sky130_fd_sc_hd__dfxtp_1
X_4923_ _4927_/A vssd1 vssd1 vccd1 vccd1 _4944_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3202__A _6024_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4854_ _5403_/B vssd1 vssd1 vccd1 vccd1 _4854_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3805_ _3803_/X _3493_/X _4402_/A vssd1 vssd1 vccd1 vccd1 _3806_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4785_ _6058_/Q _4757_/X _4767_/X _4784_/X vssd1 vssd1 vccd1 vccd1 _4785_/X sky130_fd_sc_hd__a211o_1
XFILLER_20_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3736_ _3750_/A _3736_/B vssd1 vssd1 vccd1 vccd1 _3737_/A sky130_fd_sc_hd__and2_1
X_3667_ _3667_/A vssd1 vssd1 vccd1 vccd1 _5677_/D sky130_fd_sc_hd__clkbuf_1
X_3598_ _3598_/A vssd1 vssd1 vccd1 vccd1 _3598_/X sky130_fd_sc_hd__clkbuf_2
X_5406_ _5424_/B vssd1 vssd1 vccd1 vccd1 _5417_/B sky130_fd_sc_hd__clkbuf_1
X_5337_ _6015_/Q _5336_/X _5337_/S vssd1 vssd1 vccd1 vccd1 _5338_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5268_ _5287_/C _5268_/B vssd1 vssd1 vccd1 vccd1 _5287_/D sky130_fd_sc_hd__nor2_1
XFILLER_87_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4219_ _4316_/A _5244_/B vssd1 vssd1 vccd1 vccd1 _5255_/B sky130_fd_sc_hd__or2_1
XANTENNA__4268__A2 _3459_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5199_ _5204_/A _5199_/B vssd1 vssd1 vccd1 vccd1 _5200_/A sky130_fd_sc_hd__and2_1
XFILLER_83_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_3_wb_clk_i_A _5813_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5502__A _6068_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4570_ _3139_/Y _4568_/X _4569_/Y vssd1 vssd1 vccd1 vccd1 _4575_/B sky130_fd_sc_hd__a21oi_1
X_3521_ _3346_/X _3513_/B _3342_/X vssd1 vssd1 vccd1 vccd1 _3522_/C sky130_fd_sc_hd__a21o_1
X_3452_ _3452_/A _3452_/B _3451_/X vssd1 vssd1 vccd1 vccd1 _3452_/X sky130_fd_sc_hd__or3b_1
X_3383_ _4383_/A vssd1 vssd1 vccd1 vccd1 _4366_/A sky130_fd_sc_hd__clkbuf_4
X_5122_ _5970_/Q _5122_/B vssd1 vssd1 vccd1 vccd1 _5122_/X sky130_fd_sc_hd__or2_1
XFILLER_69_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5447__A1 _5373_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5053_ _5076_/B vssd1 vssd1 vccd1 vccd1 _5066_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_84_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4004_ _5240_/A _4003_/X _4001_/Y vssd1 vssd1 vccd1 vccd1 _4452_/S sky130_fd_sc_hd__o21a_1
XFILLER_1_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5955_ _5959_/CLK _5955_/D vssd1 vssd1 vccd1 vccd1 _5955_/Q sky130_fd_sc_hd__dfxtp_1
X_4906_ _6003_/Q _5995_/Q _4914_/S vssd1 vssd1 vccd1 vccd1 _4906_/X sky130_fd_sc_hd__mux2_1
X_5886_ _6031_/CLK _5886_/D vssd1 vssd1 vccd1 vccd1 _5886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4837_ _6039_/Q _4803_/X _4804_/X vssd1 vssd1 vccd1 vccd1 _4837_/X sky130_fd_sc_hd__o21a_1
X_4768_ _4870_/A vssd1 vssd1 vccd1 vccd1 _4768_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3719_ input7/X _5691_/Q _3722_/S vssd1 vssd1 vccd1 vccd1 _3719_/X sky130_fd_sc_hd__mux2_1
X_4699_ _6098_/Q _4698_/X _4720_/S vssd1 vssd1 vccd1 vccd1 _4699_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_407 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5438__A1 _5360_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_476 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4401__A _5258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3137__C1 _3999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3152__A2 _5284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3455__A3 _3466_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4404__A2 _5254_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5740_ _6121_/CLK _5740_/D vssd1 vssd1 vccd1 vccd1 _5740_/Q sky130_fd_sc_hd__dfxtp_1
X_2952_ _5813_/Q vssd1 vssd1 vccd1 vccd1 _3296_/A sky130_fd_sc_hd__inv_2
XFILLER_22_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2883_ _3035_/C vssd1 vssd1 vccd1 vccd1 _3304_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5671_ _6091_/CLK _5671_/D vssd1 vssd1 vccd1 vccd1 _5671_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4622_ _6042_/Q _4584_/X _4610_/X _4621_/X vssd1 vssd1 vccd1 vccd1 _4622_/X sky130_fd_sc_hd__a211o_1
X_4553_ _3454_/X _3326_/A _4322_/B _4466_/X _4552_/X vssd1 vssd1 vccd1 vccd1 _4553_/X
+ sky130_fd_sc_hd__a41o_1
X_4484_ _4545_/B _4541_/A vssd1 vssd1 vccd1 vccd1 _4487_/B sky130_fd_sc_hd__nand2_1
X_3504_ _3493_/X _3410_/X _3502_/X _3503_/X vssd1 vssd1 vccd1 vccd1 _3504_/X sky130_fd_sc_hd__a211o_1
XANTENNA__5407__A _6033_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3435_ _3435_/A _5304_/A _3291_/B vssd1 vssd1 vccd1 vccd1 _3435_/X sky130_fd_sc_hd__or3b_1
XFILLER_85_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3366_ _5714_/Q vssd1 vssd1 vccd1 vccd1 _3494_/A sky130_fd_sc_hd__inv_2
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3297_ _3317_/A _3297_/B vssd1 vssd1 vccd1 vccd1 _3829_/D sky130_fd_sc_hd__or2_1
X_6085_ _6085_/CLK _6085_/D vssd1 vssd1 vccd1 vccd1 _6085_/Q sky130_fd_sc_hd__dfxtp_1
X_5105_ _5537_/B _5150_/B vssd1 vssd1 vccd1 vccd1 _5122_/B sky130_fd_sc_hd__nor2_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5036_ _5943_/Q _5942_/Q _5036_/C vssd1 vssd1 vccd1 vccd1 _5038_/A sky130_fd_sc_hd__and3_1
XFILLER_38_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5938_ _5944_/CLK _5938_/D vssd1 vssd1 vccd1 vccd1 _5938_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5869_ _5926_/CLK _5869_/D vssd1 vssd1 vccd1 vccd1 _5869_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4159__A1 _3480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput67 _5894_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[81] sky130_fd_sc_hd__buf_2
XFILLER_0_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput56 _5883_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[70] sky130_fd_sc_hd__buf_2
Xoutput78 _5905_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[92] sky130_fd_sc_hd__buf_2
XFILLER_0_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_535 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5052__A _5624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5292__C1 _4113_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input16_A la_data_in[42] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5044__C1 _5043_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3954__B _3954_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3358__C1 _3256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4131__A _4182_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3220_ _5544_/A vssd1 vssd1 vccd1 vccd1 _5638_/A sky130_fd_sc_hd__clkbuf_2
X_3151_ _3408_/B _4487_/A vssd1 vssd1 vccd1 vccd1 _4462_/S sky130_fd_sc_hd__or2_1
XFILLER_67_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_3_3__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_6_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_11_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3082_ _3480_/A _3266_/A vssd1 vssd1 vccd1 vccd1 _3082_/Y sky130_fd_sc_hd__nor2_1
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_487 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3984_ _5731_/Q _3941_/A _3953_/X _3983_/Y vssd1 vssd1 vccd1 vccd1 _3984_/X sky130_fd_sc_hd__o211a_1
XANTENNA__3210__A _6019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3597__C1 _3585_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5723_ _5736_/CLK _5723_/D vssd1 vssd1 vccd1 vccd1 _5723_/Q sky130_fd_sc_hd__dfxtp_1
X_2935_ _2949_/C _2949_/D _3312_/C _3312_/D vssd1 vssd1 vccd1 vccd1 _3317_/A sky130_fd_sc_hd__or4bb_2
X_2866_ _3298_/D vssd1 vssd1 vccd1 vccd1 _3842_/A sky130_fd_sc_hd__clkbuf_2
X_5654_ _6138_/Q _5654_/B vssd1 vssd1 vccd1 vccd1 _5654_/X sky130_fd_sc_hd__or2_1
XFILLER_30_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4605_ _5345_/A vssd1 vssd1 vccd1 vccd1 _5379_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_7_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5585_ _6098_/Q _5592_/B vssd1 vssd1 vccd1 vccd1 _5585_/X sky130_fd_sc_hd__or2_1
X_4536_ _4970_/A _4536_/B _4536_/C vssd1 vssd1 vccd1 vccd1 _4537_/A sky130_fd_sc_hd__and3_1
XFILLER_89_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4467_ _3466_/A _3483_/B _4322_/B _4466_/X _5803_/Q vssd1 vssd1 vccd1 vccd1 _4467_/X
+ sky130_fd_sc_hd__a41o_1
X_3418_ _3218_/X _3244_/C _3417_/Y vssd1 vssd1 vccd1 vccd1 _3418_/Y sky130_fd_sc_hd__a21oi_1
X_4398_ _4398_/A vssd1 vssd1 vccd1 vccd1 _5835_/D sky130_fd_sc_hd__clkbuf_1
X_3349_ _3415_/A _3854_/A _3349_/C vssd1 vssd1 vccd1 vccd1 _3349_/X sky130_fd_sc_hd__and3_1
XFILLER_58_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input8_A la_data_in[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6137_ _6138_/CLK _6137_/D vssd1 vssd1 vccd1 vccd1 _6137_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6068_ _6091_/CLK _6068_/D vssd1 vssd1 vccd1 vccd1 _6068_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_73_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5019_ _5019_/A vssd1 vssd1 vccd1 vccd1 _5937_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5329__B1 _3547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4001__B1 _4288_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3815__B1 _3525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2853__B _3518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5370_ _6023_/Q _5374_/B vssd1 vssd1 vccd1 vccd1 _5370_/X sky130_fd_sc_hd__or2_1
X_4321_ _3898_/A _3494_/B _4321_/S vssd1 vssd1 vccd1 vccd1 _4321_/X sky130_fd_sc_hd__mux2_1
X_4252_ _3873_/B _3842_/A _3315_/B vssd1 vssd1 vccd1 vccd1 _4252_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_4_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3203_ _6024_/Q _5943_/Q vssd1 vssd1 vccd1 vccd1 _3203_/X sky130_fd_sc_hd__and2_1
XFILLER_67_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3205__A _6022_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4183_ _5947_/Q _3454_/X _4196_/S vssd1 vssd1 vccd1 vccd1 _4183_/X sky130_fd_sc_hd__mux2_1
X_3134_ _4548_/A _4545_/A _3134_/C vssd1 vssd1 vccd1 vccd1 _3135_/C sky130_fd_sc_hd__nor3_1
XFILLER_82_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4059__A0 _5761_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3065_ _5277_/B _5277_/C vssd1 vssd1 vccd1 vccd1 _3066_/B sky130_fd_sc_hd__and2b_1
XANTENNA__5420__A _5461_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3967_ _3967_/A vssd1 vssd1 vccd1 vccd1 _5727_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2918_ _6012_/Q _5309_/A _6010_/Q vssd1 vssd1 vccd1 vccd1 _5323_/B sky130_fd_sc_hd__nand3b_2
X_5706_ _6085_/CLK _5706_/D vssd1 vssd1 vccd1 vccd1 _5706_/Q sky130_fd_sc_hd__dfxtp_1
X_3898_ _3898_/A _3898_/B vssd1 vssd1 vccd1 vccd1 _3903_/C sky130_fd_sc_hd__nor2_1
X_2849_ _3038_/A _5736_/Q vssd1 vssd1 vccd1 vccd1 _3118_/B sky130_fd_sc_hd__or2_1
X_5637_ _6118_/Q _5642_/B vssd1 vssd1 vccd1 vccd1 _5637_/X sky130_fd_sc_hd__or2_1
X_5568_ _6092_/Q _5570_/B vssd1 vssd1 vccd1 vccd1 _5568_/X sky130_fd_sc_hd__or2_1
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4519_ _4504_/Y _4517_/X _4518_/Y _4511_/A _5863_/Q vssd1 vssd1 vccd1 vccd1 _4520_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_2_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_37_wb_clk_i_A clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_5499_ _5353_/X _5493_/X _5498_/X _5488_/X vssd1 vssd1 vccd1 vccd1 _6066_/D sky130_fd_sc_hd__o211a_1
XFILLER_77_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3115__A _5736_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4645__S _4645_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3935__D _6121_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3500__A2 _3411_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5253__A2 _5278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4870_ _4870_/A vssd1 vssd1 vccd1 vccd1 _4870_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3821_ _3821_/A _3891_/B _3821_/C vssd1 vssd1 vccd1 vccd1 _3821_/X sky130_fd_sc_hd__and3_1
XFILLER_20_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3752_ _3770_/A vssd1 vssd1 vccd1 vccd1 _3768_/A sky130_fd_sc_hd__clkbuf_1
X_3683_ _3587_/A _5682_/Q _3697_/S vssd1 vssd1 vccd1 vccd1 _3684_/B sky130_fd_sc_hd__mux2_1
X_5422_ _6039_/Q _5424_/B vssd1 vssd1 vccd1 vccd1 _5422_/X sky130_fd_sc_hd__or2_1
X_5353_ input6/X vssd1 vssd1 vccd1 vccd1 _5353_/X sky130_fd_sc_hd__clkbuf_2
X_4304_ _3357_/X _3497_/X _4294_/A vssd1 vssd1 vccd1 vccd1 _4306_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__5415__A _6036_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5284_ _5284_/A _5284_/B _5284_/C vssd1 vssd1 vccd1 vccd1 _6008_/D sky130_fd_sc_hd__nor3_1
XFILLER_87_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4235_ _6132_/Q _6122_/Q _4235_/C _6128_/Q vssd1 vssd1 vccd1 vccd1 _5252_/B sky130_fd_sc_hd__or4_1
X_4166_ _5660_/Q _5791_/Q _4179_/S vssd1 vssd1 vccd1 vccd1 _4166_/X sky130_fd_sc_hd__mux2_1
X_3117_ _3117_/A _3117_/B vssd1 vssd1 vccd1 vccd1 _3117_/Y sky130_fd_sc_hd__nor2_1
XFILLER_82_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4097_ _5772_/Q _4096_/X _4097_/S vssd1 vssd1 vccd1 vccd1 _4098_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3589__B _3765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5150__A _5405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3048_ _3043_/X _3046_/Y _3047_/X vssd1 vssd1 vccd1 vccd1 _3059_/C sky130_fd_sc_hd__o21bai_1
XFILLER_63_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3558__A2 _4331_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4755__A1 _5891_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4999_ _4999_/A _4999_/B vssd1 vssd1 vccd1 vccd1 _5931_/D sky130_fd_sc_hd__nor2_1
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5468__C1 _5461_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3719__S _3722_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4746__A1 _6030_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4020_ _4020_/A vssd1 vssd1 vccd1 vccd1 _5749_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5971_ _5975_/CLK _5971_/D vssd1 vssd1 vccd1 vccd1 _5971_/Q sky130_fd_sc_hd__dfxtp_1
X_4922_ _5873_/Q _5852_/Q vssd1 vssd1 vccd1 vccd1 _4927_/A sky130_fd_sc_hd__nand2_1
X_4853_ _5971_/Q _4808_/X _4818_/X _4852_/X vssd1 vssd1 vccd1 vccd1 _4853_/X sky130_fd_sc_hd__a211o_1
X_3804_ _4432_/S _3379_/A _3525_/A vssd1 vssd1 vccd1 vccd1 _4402_/A sky130_fd_sc_hd__o21ai_1
X_4784_ _4768_/X _4782_/X _4783_/X _4773_/X vssd1 vssd1 vccd1 vccd1 _4784_/X sky130_fd_sc_hd__o211a_1
X_3735_ _5373_/A _5696_/Q _3735_/S vssd1 vssd1 vccd1 vccd1 _3736_/B sky130_fd_sc_hd__mux2_1
X_3666_ _3666_/A _3666_/B vssd1 vssd1 vccd1 vccd1 _3667_/A sky130_fd_sc_hd__and2_1
X_5405_ _5603_/A _5405_/B vssd1 vssd1 vccd1 vccd1 _5424_/B sky130_fd_sc_hd__nor2_1
X_3597_ _3587_/X _3592_/X _3596_/X _3585_/X vssd1 vssd1 vccd1 vccd1 _5658_/D sky130_fd_sc_hd__o211a_1
XFILLER_87_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5336_ _6067_/Q _6014_/Q _5336_/S vssd1 vssd1 vccd1 vccd1 _5336_/X sky130_fd_sc_hd__mux2_1
X_5267_ _5339_/S _3067_/A _5287_/A vssd1 vssd1 vccd1 vccd1 _5278_/D sky130_fd_sc_hd__a21o_1
XFILLER_87_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4218_ _4218_/A _4218_/B vssd1 vssd1 vccd1 vccd1 _5244_/B sky130_fd_sc_hd__nand2_2
X_5198_ _5075_/A _5996_/Q _5198_/S vssd1 vssd1 vccd1 vccd1 _5199_/B sky130_fd_sc_hd__mux2_1
XFILLER_68_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4149_ _6137_/Q _5786_/Q _4162_/S vssd1 vssd1 vccd1 vccd1 _4149_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5153__A1 _5045_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input46_A wbs_sel_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_471 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_40 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5392__A1 _5389_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3520_ _3520_/A _3520_/B vssd1 vssd1 vccd1 vccd1 _3520_/X sky130_fd_sc_hd__or2_1
XFILLER_6_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3451_ _3460_/A _5320_/A _3460_/C _3451_/D vssd1 vssd1 vccd1 vccd1 _3451_/X sky130_fd_sc_hd__or4_1
X_3382_ _5257_/A vssd1 vssd1 vccd1 vccd1 _4383_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_41_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5121_ _5072_/X _5104_/A _5120_/X _5114_/X vssd1 vssd1 vccd1 vccd1 _5969_/D sky130_fd_sc_hd__o211a_1
XFILLER_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5052_ _5624_/A _5150_/B vssd1 vssd1 vccd1 vccd1 _5076_/B sky130_fd_sc_hd__nor2_1
X_4003_ _4236_/A _4003_/B vssd1 vssd1 vccd1 vccd1 _4003_/X sky130_fd_sc_hd__or2_1
XFILLER_92_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5954_ _6064_/CLK _5954_/D vssd1 vssd1 vccd1 vccd1 _5954_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_52_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4905_ _5906_/Q _4858_/X _4903_/X _4904_/X vssd1 vssd1 vccd1 vccd1 _5906_/D sky130_fd_sc_hd__a22o_1
X_5885_ _6031_/CLK _5885_/D vssd1 vssd1 vccd1 vccd1 _5885_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4044__A _4095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4836_ _6063_/Q _4808_/X _4818_/X _4835_/X vssd1 vssd1 vccd1 vccd1 _4836_/X sky130_fd_sc_hd__a211o_1
X_4767_ _4869_/A vssd1 vssd1 vccd1 vccd1 _4767_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3718_ _5171_/A _3718_/B vssd1 vssd1 vccd1 vccd1 _5690_/D sky130_fd_sc_hd__nor2_1
XFILLER_20_14 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4698_ _6134_/Q _4697_/X _4719_/S vssd1 vssd1 vccd1 vccd1 _4698_/X sky130_fd_sc_hd__mux2_1
X_3649_ _3649_/A vssd1 vssd1 vccd1 vccd1 _5672_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5319_ _4231_/A _3322_/X _3439_/A _4464_/X vssd1 vssd1 vccd1 vccd1 _5320_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2962__A _2994_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3909__C1 _4554_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_3_2__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5813_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__5513__A _5579_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3968__A _5188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2951_ _3850_/C vssd1 vssd1 vccd1 vccd1 _5327_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_34_179 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5670_ _6091_/CLK _5670_/D vssd1 vssd1 vccd1 vccd1 _5670_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_32_wb_clk_i _5836_/CLK vssd1 vssd1 vccd1 vccd1 _6109_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_89_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2882_ _3853_/C _3833_/C _3256_/A vssd1 vssd1 vccd1 vccd1 _3035_/C sky130_fd_sc_hd__and3_1
X_4621_ _4611_/X _4615_/X _4618_/X _4620_/X vssd1 vssd1 vccd1 vccd1 _4621_/X sky130_fd_sc_hd__o211a_1
XANTENNA__5365__A1 _5363_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4552_ _4551_/X _5796_/Q vssd1 vssd1 vccd1 vccd1 _4552_/X sky130_fd_sc_hd__and2b_1
X_4483_ _4481_/X _4482_/X _3245_/X vssd1 vssd1 vccd1 vccd1 _5857_/D sky130_fd_sc_hd__o21a_1
X_3503_ _3494_/A _3274_/C _3891_/B _3269_/X vssd1 vssd1 vccd1 vccd1 _3503_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3853__D _3897_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3434_ _3434_/A vssd1 vssd1 vccd1 vccd1 _3434_/Y sky130_fd_sc_hd__inv_2
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3365_ _4432_/S vssd1 vssd1 vccd1 vccd1 _4409_/S sky130_fd_sc_hd__clkbuf_2
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3296_ _3296_/A _3296_/B vssd1 vssd1 vccd1 vccd1 _4283_/B sky130_fd_sc_hd__nand2_1
X_6084_ _6087_/CLK _6084_/D vssd1 vssd1 vccd1 vccd1 _6084_/Q sky130_fd_sc_hd__dfxtp_1
X_5104_ _5104_/A vssd1 vssd1 vccd1 vccd1 _5104_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5035_ _5035_/A _5035_/B vssd1 vssd1 vccd1 vccd1 _5942_/D sky130_fd_sc_hd__nor2_1
XFILLER_57_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5937_ _5945_/CLK _5937_/D vssd1 vssd1 vccd1 vccd1 _5937_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5868_ _5926_/CLK _5868_/D vssd1 vssd1 vccd1 vccd1 _5868_/Q sky130_fd_sc_hd__dfxtp_1
X_4819_ _4870_/A vssd1 vssd1 vccd1 vccd1 _4819_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__5356__A1 _5353_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5799_ _5959_/CLK _5799_/D vssd1 vssd1 vccd1 vccd1 _5799_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4564__C1 _3723_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5108__A1 _5045_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput57 _5884_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[71] sky130_fd_sc_hd__buf_2
XFILLER_0_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput68 _5895_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[82] sky130_fd_sc_hd__buf_2
Xoutput79 _5906_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[93] sky130_fd_sc_hd__buf_2
XFILLER_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5595__A1 _5396_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2867__A _3842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3150_ _3391_/A _5743_/Q vssd1 vssd1 vccd1 vccd1 _4487_/A sky130_fd_sc_hd__nand2_1
XFILLER_67_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3081_ _3480_/A _3081_/B vssd1 vssd1 vccd1 vccd1 _3081_/X sky130_fd_sc_hd__and2_1
XFILLER_54_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4086__A1 _3287_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3983_ _5731_/Q _3983_/B vssd1 vssd1 vccd1 vccd1 _3983_/Y sky130_fd_sc_hd__nand2_1
X_5722_ _5736_/CLK _5722_/D vssd1 vssd1 vccd1 vccd1 _5722_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2934_ _5814_/Q vssd1 vssd1 vccd1 vccd1 _3312_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_50_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2865_ _5808_/Q _5807_/Q _5806_/Q _4249_/B vssd1 vssd1 vccd1 vccd1 _3298_/D sky130_fd_sc_hd__and4bb_1
X_5653_ _5393_/X _3576_/A _5652_/X _5172_/X vssd1 vssd1 vccd1 vccd1 _6137_/D sky130_fd_sc_hd__o211a_1
X_4604_ _4604_/A _4604_/B vssd1 vssd1 vccd1 vccd1 _5345_/A sky130_fd_sc_hd__or2_1
X_5584_ _5376_/X _5580_/X _5583_/X _5571_/X vssd1 vssd1 vccd1 vccd1 _6097_/D sky130_fd_sc_hd__o211a_1
XFILLER_30_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4535_ _4535_/A _4541_/B vssd1 vssd1 vccd1 vccd1 _4536_/C sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_27_wb_clk_i_A clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xuser_proj_example_190 vssd1 vssd1 vccd1 vccd1 user_proj_example_190/HI la_data_out[97]
+ sky130_fd_sc_hd__conb_1
X_4466_ _4466_/A _4466_/B _4466_/C vssd1 vssd1 vccd1 vccd1 _4466_/X sky130_fd_sc_hd__and3_1
X_3417_ _4982_/B vssd1 vssd1 vccd1 vccd1 _3417_/Y sky130_fd_sc_hd__inv_2
X_4397_ _5835_/Q _4396_/X _4397_/S vssd1 vssd1 vccd1 vccd1 _4398_/A sky130_fd_sc_hd__mux2_1
X_3348_ _5240_/A _3814_/C _3340_/X _3347_/X vssd1 vssd1 vccd1 vccd1 _3348_/X sky130_fd_sc_hd__a211o_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6136_ _6138_/CLK _6136_/D vssd1 vssd1 vccd1 vccd1 _6136_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3279_ _4233_/A _3274_/X _3277_/Y _3415_/A vssd1 vssd1 vccd1 vccd1 _3279_/X sky130_fd_sc_hd__a2bb2o_1
X_6067_ _6067_/CLK _6067_/D vssd1 vssd1 vccd1 vccd1 _6067_/Q sky130_fd_sc_hd__dfxtp_2
X_5018_ _5023_/C _5025_/B _5018_/C vssd1 vssd1 vccd1 vccd1 _5019_/A sky130_fd_sc_hd__and3b_1
XFILLER_26_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5047__B _5201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4304__A2 _3497_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5501__A1 _5357_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3512__B1 _3245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_514 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3311__A _4438_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4320_ _3275_/X _3079_/B _3276_/Y vssd1 vssd1 vccd1 vccd1 _4320_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_4_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4251_ _4251_/A vssd1 vssd1 vccd1 vccd1 _4970_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_86_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3503__B1 _3269_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3202_ _6024_/Q _5943_/Q vssd1 vssd1 vccd1 vccd1 _3202_/Y sky130_fd_sc_hd__nor2_1
XFILLER_67_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4182_ _4182_/A vssd1 vssd1 vccd1 vccd1 _4196_/S sky130_fd_sc_hd__clkbuf_2
X_3133_ _5868_/Q _5867_/Q _5865_/Q _5866_/Q vssd1 vssd1 vccd1 vccd1 _3134_/C sky130_fd_sc_hd__or4b_1
X_3064_ _6007_/Q vssd1 vssd1 vccd1 vccd1 _5277_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_70_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3221__A _5638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3966_ _3966_/A _3966_/B vssd1 vssd1 vccd1 vccd1 _3967_/A sky130_fd_sc_hd__and2_1
X_2917_ _2917_/A vssd1 vssd1 vccd1 vccd1 _3460_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5705_ _5892_/CLK _5705_/D vssd1 vssd1 vccd1 vccd1 _5705_/Q sky130_fd_sc_hd__dfxtp_1
X_3897_ _3897_/A _3897_/B _4259_/A _3897_/D vssd1 vssd1 vccd1 vccd1 _3898_/B sky130_fd_sc_hd__or4_1
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5148__A _5405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5636_ _5363_/X _5623_/X _5635_/X _5627_/X vssd1 vssd1 vccd1 vccd1 _6117_/D sky130_fd_sc_hd__o211a_1
X_2848_ _5848_/Q vssd1 vssd1 vccd1 vccd1 _3038_/A sky130_fd_sc_hd__buf_2
X_5567_ _5357_/X _5559_/X _5566_/X _5556_/X vssd1 vssd1 vccd1 vccd1 _6091_/D sky130_fd_sc_hd__o211a_1
X_4518_ _5863_/Q _5862_/Q _4518_/C _4518_/D vssd1 vssd1 vccd1 vccd1 _4518_/Y sky130_fd_sc_hd__nand4_1
X_5498_ _6066_/Q _5505_/B vssd1 vssd1 vccd1 vccd1 _5498_/X sky130_fd_sc_hd__or2_1
X_4449_ _3820_/A _3331_/X _4443_/X _4448_/X vssd1 vssd1 vccd1 vccd1 _4449_/X sky130_fd_sc_hd__a31o_1
XFILLER_58_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6119_ _6135_/CLK _6119_/D vssd1 vssd1 vccd1 vccd1 _6119_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2954__B _3836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4446__D1 _4466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4213__A1 _3037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3820_ _3820_/A _3820_/B _4229_/A vssd1 vssd1 vccd1 vccd1 _3820_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__2880__A _2880_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3751_ _3751_/A vssd1 vssd1 vccd1 vccd1 _5700_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4764__A2 _4757_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3682_ _3707_/S vssd1 vssd1 vccd1 vccd1 _3697_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_3_2__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5421_ _3611_/X _5404_/A _5419_/X _5420_/X vssd1 vssd1 vccd1 vccd1 _6038_/D sky130_fd_sc_hd__o211a_1
X_5352_ _5342_/X _5347_/X _5351_/X _5169_/X vssd1 vssd1 vccd1 vccd1 _6017_/D sky130_fd_sc_hd__o211a_1
X_4303_ _3405_/A _3497_/X _4233_/C vssd1 vssd1 vccd1 vccd1 _4306_/B sky130_fd_sc_hd__a21oi_1
X_5283_ _5297_/C _5278_/Y _5282_/X _5262_/X vssd1 vssd1 vccd1 vccd1 _5284_/C sky130_fd_sc_hd__o211a_1
X_4234_ _5256_/B _4234_/B vssd1 vssd1 vccd1 vccd1 _4243_/A sky130_fd_sc_hd__and2_1
X_4165_ _4182_/A vssd1 vssd1 vccd1 vccd1 _4179_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_82_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3116_ _3116_/A vssd1 vssd1 vccd1 vccd1 _3117_/B sky130_fd_sc_hd__clkbuf_2
X_4096_ _5958_/Q _5771_/Q _4110_/S vssd1 vssd1 vccd1 vccd1 _4096_/X sky130_fd_sc_hd__mux2_1
X_3047_ _3047_/A vssd1 vssd1 vccd1 vccd1 _3047_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4452__A1 _4449_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4998_ _5931_/Q _5000_/C _4990_/X vssd1 vssd1 vccd1 vccd1 _4999_/B sky130_fd_sc_hd__o21ai_1
X_3949_ _5724_/Q _3932_/A _3945_/X _5723_/Q vssd1 vssd1 vccd1 vccd1 _3950_/B sky130_fd_sc_hd__a22o_1
XFILLER_23_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5619_ _3614_/X _5602_/A _5618_/X _5612_/X vssd1 vssd1 vccd1 vccd1 _6111_/D sky130_fd_sc_hd__o211a_1
XFILLER_2_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_520 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_57_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6077_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_84_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5970_ _5975_/CLK _5970_/D vssd1 vssd1 vccd1 vccd1 _5970_/Q sky130_fd_sc_hd__dfxtp_1
X_4921_ _5908_/Q _4623_/X _4919_/X _4920_/X vssd1 vssd1 vccd1 vccd1 _5908_/D sky130_fd_sc_hd__a22o_1
X_4852_ _4819_/X _4850_/X _4851_/X _4824_/X vssd1 vssd1 vccd1 vccd1 _4852_/X sky130_fd_sc_hd__o211a_1
XFILLER_60_383 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3803_ _4409_/S _3800_/Y _3801_/X _3802_/X vssd1 vssd1 vccd1 vccd1 _3803_/X sky130_fd_sc_hd__a31o_1
X_4783_ _6082_/Q _4783_/B vssd1 vssd1 vccd1 vccd1 _4783_/X sky130_fd_sc_hd__or2_1
XFILLER_9_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3734_ _3770_/A vssd1 vssd1 vccd1 vccd1 _3750_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_9_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3665_ _5389_/A _5677_/Q _3669_/S vssd1 vssd1 vccd1 vccd1 _3666_/B sky130_fd_sc_hd__mux2_1
XANTENNA__5426__A _5471_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5404_ _5404_/A vssd1 vssd1 vccd1 vccd1 _5404_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3596_ _5658_/Q _3608_/B vssd1 vssd1 vccd1 vccd1 _3596_/X sky130_fd_sc_hd__or2_1
X_5335_ _5335_/A vssd1 vssd1 vccd1 vccd1 _6014_/D sky130_fd_sc_hd__clkbuf_1
X_5266_ _5294_/S vssd1 vssd1 vccd1 vccd1 _5266_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4217_ _4217_/A _4217_/B vssd1 vssd1 vccd1 vccd1 _4316_/A sky130_fd_sc_hd__nand2_1
X_5197_ _5197_/A vssd1 vssd1 vccd1 vccd1 _5995_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4148_ _4182_/A vssd1 vssd1 vccd1 vccd1 _4162_/S sky130_fd_sc_hd__buf_2
X_4079_ _6110_/Q _5766_/Q _4092_/S vssd1 vssd1 vccd1 vccd1 _4079_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_1__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_5_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_input39_A la_data_in[63] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3450_ _3447_/X _3449_/X _2955_/X vssd1 vssd1 vccd1 vccd1 _3452_/B sky130_fd_sc_hd__o21a_1
XFILLER_6_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3381_ _4235_/C vssd1 vssd1 vccd1 vccd1 _5257_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5120_ _5969_/Q _5122_/B vssd1 vssd1 vccd1 vccd1 _5120_/X sky130_fd_sc_hd__or2_1
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5051_ _5051_/A vssd1 vssd1 vccd1 vccd1 _5150_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4002_ _4002_/A _6124_/Q _6127_/Q _6128_/Q vssd1 vssd1 vccd1 vccd1 _4003_/B sky130_fd_sc_hd__or4_1
XFILLER_77_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5953_ _6064_/CLK _5953_/D vssd1 vssd1 vccd1 vccd1 _5953_/Q sky130_fd_sc_hd__dfxtp_1
X_4904_ _5984_/Q _5379_/B _4607_/A vssd1 vssd1 vccd1 vccd1 _4904_/X sky130_fd_sc_hd__o21a_1
XFILLER_21_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5884_ _6027_/CLK _5884_/D vssd1 vssd1 vccd1 vccd1 _5884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4835_ _4819_/X _4833_/X _4834_/X _4824_/X vssd1 vssd1 vccd1 vccd1 _4835_/X sky130_fd_sc_hd__o211a_1
XFILLER_21_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4766_ _5892_/Q _4756_/X _4764_/X _4765_/Y vssd1 vssd1 vccd1 vccd1 _5892_/D sky130_fd_sc_hd__a22o_1
X_3717_ _4575_/A _3716_/X _5875_/Q vssd1 vssd1 vccd1 vccd1 _3718_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__5156__A _5981_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4697_ _5698_/Q _5675_/Q _4697_/S vssd1 vssd1 vccd1 vccd1 _4697_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3648_ _3648_/A _3648_/B vssd1 vssd1 vccd1 vccd1 _3649_/A sky130_fd_sc_hd__and2_1
XANTENNA__5540__C1 _5529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3579_ _5654_/B vssd1 vssd1 vccd1 vccd1 _5648_/B sky130_fd_sc_hd__clkbuf_1
X_5318_ _5315_/A _5266_/X _5317_/Y _5169_/X vssd1 vssd1 vccd1 vccd1 _6011_/D sky130_fd_sc_hd__o211a_1
XFILLER_88_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5603__B _5603_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5249_ _5249_/A _5258_/B _5269_/C vssd1 vssd1 vccd1 vccd1 _5278_/C sky130_fd_sc_hd__or3_1
XANTENNA__3404__A _3842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_2_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6117_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_16_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3606__C1 _3585_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3385__A1 _4409_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5513__B _5535_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_423 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5598__C1 _5597_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2950_ _2950_/A _2950_/B _3312_/B _3312_/C vssd1 vssd1 vccd1 vccd1 _3850_/C sky130_fd_sc_hd__or4b_2
XFILLER_62_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2881_ _3838_/A _3836_/A vssd1 vssd1 vccd1 vccd1 _3256_/A sky130_fd_sc_hd__nor2_2
XFILLER_15_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4620_ _4824_/A vssd1 vssd1 vccd1 vccd1 _4620_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4551_ _3483_/B _3482_/Y _4550_/Y _4464_/X _4466_/X vssd1 vssd1 vccd1 vccd1 _4551_/X
+ sky130_fd_sc_hd__o221a_1
X_4482_ _4480_/A _3561_/A _3135_/X vssd1 vssd1 vccd1 vccd1 _4482_/X sky130_fd_sc_hd__o21a_1
X_3502_ _3502_/A _3502_/B vssd1 vssd1 vccd1 vccd1 _3502_/X sky130_fd_sc_hd__and2_1
X_3433_ _3431_/X _3432_/X _3046_/A vssd1 vssd1 vccd1 vccd1 _3433_/Y sky130_fd_sc_hd__a21oi_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3364_ _5258_/A vssd1 vssd1 vccd1 vccd1 _4432_/S sky130_fd_sc_hd__clkbuf_2
X_5103_ _5535_/B _5148_/B vssd1 vssd1 vccd1 vccd1 _5104_/A sky130_fd_sc_hd__or2_1
XFILLER_85_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3295_ _5241_/C _5247_/B _3350_/B _2972_/X vssd1 vssd1 vccd1 vccd1 _3300_/C sky130_fd_sc_hd__a31o_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6083_ _6085_/CLK _6083_/D vssd1 vssd1 vccd1 vccd1 _6083_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5034_ _5942_/Q _5036_/C _5020_/X vssd1 vssd1 vccd1 vccd1 _5035_/B sky130_fd_sc_hd__o21ai_1
XFILLER_80_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5936_ _5945_/CLK _5936_/D vssd1 vssd1 vccd1 vccd1 _5936_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_56_wb_clk_i_A clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_5867_ _5926_/CLK _5867_/D vssd1 vssd1 vccd1 vccd1 _5867_/Q sky130_fd_sc_hd__dfxtp_1
X_5798_ _5959_/CLK _5798_/D vssd1 vssd1 vccd1 vccd1 _5798_/Q sky130_fd_sc_hd__dfxtp_1
X_4818_ _4869_/A vssd1 vssd1 vccd1 vccd1 _4818_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4749_ _5656_/Q _4748_/X _4770_/S vssd1 vssd1 vccd1 vccd1 _4749_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput58 _5885_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[72] sky130_fd_sc_hd__buf_2
XANTENNA__4867__A1 _5980_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput69 _5896_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[83] sky130_fd_sc_hd__buf_2
XANTENNA__5292__A1 _5327_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3080_ _5241_/A vssd1 vssd1 vccd1 vccd1 _3480_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_67_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3982_ _3982_/A vssd1 vssd1 vccd1 vccd1 _5731_/D sky130_fd_sc_hd__clkbuf_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2933_ _2933_/A _2942_/A vssd1 vssd1 vccd1 vccd1 _2936_/A sky130_fd_sc_hd__or2_1
XFILLER_62_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5721_ _5777_/CLK _5721_/D vssd1 vssd1 vccd1 vccd1 _5721_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2864_ _5805_/Q vssd1 vssd1 vccd1 vccd1 _4249_/B sky130_fd_sc_hd__clkbuf_1
X_5652_ _6137_/Q _5654_/B vssd1 vssd1 vccd1 vccd1 _5652_/X sky130_fd_sc_hd__or2_1
XANTENNA__4322__B _4322_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5583_ _6097_/Q _5592_/B vssd1 vssd1 vccd1 vccd1 _5583_/X sky130_fd_sc_hd__or2_1
X_4603_ _6041_/Q _4584_/X _4599_/X _4602_/X vssd1 vssd1 vccd1 vccd1 _4603_/X sky130_fd_sc_hd__a211o_1
X_4534_ _4534_/A _4534_/B _4534_/C vssd1 vssd1 vccd1 vccd1 _4541_/B sky130_fd_sc_hd__and3_1
XFILLER_7_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_proj_example_180 vssd1 vssd1 vccd1 vccd1 user_proj_example_180/HI la_data_out[55]
+ sky130_fd_sc_hd__conb_1
X_4465_ _3438_/A _3322_/X _4464_/X vssd1 vssd1 vccd1 vccd1 _4466_/C sky130_fd_sc_hd__a21bo_1
Xuser_proj_example_191 vssd1 vssd1 vccd1 vccd1 user_proj_example_191/HI la_data_out[98]
+ sky130_fd_sc_hd__conb_1
X_3416_ _3272_/B _3409_/X _3415_/Y vssd1 vssd1 vccd1 vccd1 _6130_/D sky130_fd_sc_hd__o21ai_1
X_4396_ _6057_/Q _5834_/Q _4396_/S vssd1 vssd1 vccd1 vccd1 _4396_/X sky130_fd_sc_hd__mux2_1
X_3347_ _3415_/A _3076_/Y _3342_/X _3346_/X vssd1 vssd1 vccd1 vccd1 _3347_/X sky130_fd_sc_hd__a211o_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6135_ _6135_/CLK _6135_/D vssd1 vssd1 vccd1 vccd1 _6135_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6066_ _6067_/CLK _6066_/D vssd1 vssd1 vccd1 vccd1 _6066_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_85_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3278_ _6130_/Q vssd1 vssd1 vccd1 vccd1 _3415_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5017_ _5936_/Q _4946_/C _4972_/A _5937_/Q vssd1 vssd1 vccd1 vccd1 _5018_/C sky130_fd_sc_hd__a31o_1
XFILLER_45_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3401__B _3802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5919_ _5920_/CLK _5919_/D vssd1 vssd1 vccd1 vccd1 _5919_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3129__A _5667_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input21_A la_data_in[47] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3815__A2 _3379_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4394__S _4397_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3039__A _3049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4250_ _4276_/A _4250_/B _4275_/C vssd1 vssd1 vccd1 vccd1 _5806_/D sky130_fd_sc_hd__nor3_1
XFILLER_79_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3201_ _6023_/Q _3198_/Y _5937_/Q _5354_/A _3200_/Y vssd1 vssd1 vccd1 vccd1 _3214_/A
+ sky130_fd_sc_hd__o221a_1
X_4181_ _4181_/A vssd1 vssd1 vccd1 vccd1 _5796_/D sky130_fd_sc_hd__clkbuf_1
X_3132_ _5869_/Q vssd1 vssd1 vccd1 vccd1 _4545_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_67_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3063_ _5297_/B _5281_/A _3063_/C vssd1 vssd1 vccd1 vccd1 _3373_/A sky130_fd_sc_hd__and3b_1
XFILLER_27_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3019__B1 _3432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3965_ _5727_/Q _3964_/X _3945_/X _5726_/Q vssd1 vssd1 vccd1 vccd1 _3966_/B sky130_fd_sc_hd__a22o_1
X_3896_ _3896_/A vssd1 vssd1 vccd1 vccd1 _4259_/A sky130_fd_sc_hd__clkbuf_2
X_2916_ _2950_/B _3312_/B _2950_/A vssd1 vssd1 vccd1 vccd1 _2917_/A sky130_fd_sc_hd__and3b_1
XANTENNA__4333__A _6068_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5704_ _5892_/CLK _5704_/D vssd1 vssd1 vccd1 vccd1 _5704_/Q sky130_fd_sc_hd__dfxtp_1
X_2847_ _3508_/B _3507_/A vssd1 vssd1 vccd1 vccd1 _2853_/C sky130_fd_sc_hd__nand2_1
XFILLER_31_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5635_ _6117_/Q _5635_/B vssd1 vssd1 vccd1 vccd1 _5635_/X sky130_fd_sc_hd__or2_1
XFILLER_12_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3891__B _3891_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5566_ _6091_/Q _5570_/B vssd1 vssd1 vccd1 vccd1 _5566_/X sky130_fd_sc_hd__or2_1
X_4517_ _5862_/Q _4518_/C _5860_/Q _5863_/Q vssd1 vssd1 vccd1 vccd1 _4517_/X sky130_fd_sc_hd__a31o_1
X_5497_ _5342_/X _5493_/X _5496_/X _5488_/X vssd1 vssd1 vccd1 vccd1 _6065_/D sky130_fd_sc_hd__o211a_1
X_4448_ _3897_/D _4443_/X _4446_/X _4447_/X vssd1 vssd1 vccd1 vccd1 _4448_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_77_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4379_ _4379_/A vssd1 vssd1 vccd1 vccd1 _5829_/D sky130_fd_sc_hd__clkbuf_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6118_ _6118_/CLK _6118_/D vssd1 vssd1 vccd1 vccd1 _6118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6049_ _6080_/CLK _6049_/D vssd1 vssd1 vccd1 vccd1 _6049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5486__A1 _3611_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3750_ _3750_/A _3750_/B vssd1 vssd1 vccd1 vccd1 _3751_/A sky130_fd_sc_hd__and2_1
XFILLER_13_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4153__A _4170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3681_ _3765_/A _5174_/A vssd1 vssd1 vccd1 vccd1 _3707_/S sky130_fd_sc_hd__nand2_1
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5420_ _5461_/A vssd1 vssd1 vccd1 vccd1 _5420_/X sky130_fd_sc_hd__clkbuf_2
X_5351_ _6017_/Q _5367_/B vssd1 vssd1 vccd1 vccd1 _5351_/X sky130_fd_sc_hd__or2_1
X_5282_ _5297_/C _5281_/B _5281_/Y _5244_/B vssd1 vssd1 vccd1 vccd1 _5282_/X sky130_fd_sc_hd__a211o_1
X_4302_ _3266_/A _3079_/B _4233_/A vssd1 vssd1 vccd1 vccd1 _4306_/A sky130_fd_sc_hd__a21oi_1
X_4233_ _4233_/A _4233_/B _4233_/C vssd1 vssd1 vccd1 vccd1 _4233_/X sky130_fd_sc_hd__and3_1
XFILLER_4_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3488__B1 _3269_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4164_ _4164_/A vssd1 vssd1 vccd1 vccd1 _5791_/D sky130_fd_sc_hd__clkbuf_1
X_3115_ _5736_/Q vssd1 vssd1 vccd1 vccd1 _3938_/A sky130_fd_sc_hd__buf_2
X_4095_ _4095_/A vssd1 vssd1 vccd1 vccd1 _4110_/S sky130_fd_sc_hd__buf_2
X_3046_ _3046_/A _3046_/B vssd1 vssd1 vccd1 vccd1 _3046_/Y sky130_fd_sc_hd__nor2_1
XFILLER_55_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3232__A _6029_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4997_ _5931_/Q _5000_/C vssd1 vssd1 vccd1 vccd1 _4999_/A sky130_fd_sc_hd__and2_1
X_3948_ _3948_/A vssd1 vssd1 vccd1 vccd1 _5723_/D sky130_fd_sc_hd__clkbuf_1
X_3879_ _3851_/C _3891_/A _4466_/A _3432_/B vssd1 vssd1 vccd1 vccd1 _3879_/Y sky130_fd_sc_hd__o211ai_1
X_5618_ _6111_/Q _5620_/B vssd1 vssd1 vccd1 vccd1 _5618_/X sky130_fd_sc_hd__or2_1
XANTENNA__4912__B1 _4607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5549_ _6085_/Q _5549_/B vssd1 vssd1 vccd1 vccd1 _5549_/X sky130_fd_sc_hd__or2_1
XFILLER_3_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_3_0__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_4_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__5468__A1 _3582_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5622__A _5622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3142__A _3723_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2981__A _3824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3651__A0 _5373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3317__A _3317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5459__A1 _5389_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_26_wb_clk_i clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5922_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_49_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output52_A _5879_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4148__A _4182_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4920_ _5986_/Q _5379_/B _4607_/A vssd1 vssd1 vccd1 vccd1 _4920_/X sky130_fd_sc_hd__o21a_1
X_4851_ _5963_/Q _4885_/B vssd1 vssd1 vccd1 vccd1 _4851_/X sky130_fd_sc_hd__or2_1
X_3802_ _5976_/Q _3802_/B vssd1 vssd1 vccd1 vccd1 _3802_/X sky130_fd_sc_hd__and2_1
XFILLER_60_395 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4782_ _6106_/Q _4780_/X _4822_/S vssd1 vssd1 vccd1 vccd1 _4782_/X sky130_fd_sc_hd__mux2_1
X_3733_ _3733_/A vssd1 vssd1 vccd1 vccd1 _5695_/D sky130_fd_sc_hd__clkbuf_1
X_3664_ _3664_/A vssd1 vssd1 vccd1 vccd1 _5676_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4611__A _4717_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5403_ _5601_/A _5403_/B vssd1 vssd1 vccd1 vccd1 _5404_/A sky130_fd_sc_hd__or2_1
X_3595_ _3618_/B vssd1 vssd1 vccd1 vccd1 _3608_/B sky130_fd_sc_hd__clkbuf_1
X_5334_ _6014_/Q _5333_/X _5337_/S vssd1 vssd1 vccd1 vccd1 _5335_/A sky130_fd_sc_hd__mux2_1
X_5265_ _5243_/A _5263_/X _5264_/X vssd1 vssd1 vccd1 vccd1 _6006_/D sky130_fd_sc_hd__o21ba_1
XFILLER_87_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4216_ _3901_/B _4215_/X _4287_/A vssd1 vssd1 vccd1 vccd1 _4227_/B sky130_fd_sc_hd__o21ai_1
X_5196_ _5204_/A _5196_/B vssd1 vssd1 vccd1 vccd1 _5197_/A sky130_fd_sc_hd__and2_1
XFILLER_68_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4147_ _4147_/A vssd1 vssd1 vccd1 vccd1 _5786_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3897__A _3897_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4078_ _4095_/A vssd1 vssd1 vccd1 vccd1 _4092_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_70_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3029_ _3826_/C vssd1 vssd1 vccd1 vccd1 _3264_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_43_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3397__C1 _3117_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5613__A1 _3604_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3380_ _5234_/A _3380_/B _3518_/B vssd1 vssd1 vccd1 vccd1 _3380_/Y sky130_fd_sc_hd__nor3_1
XFILLER_69_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5050_ _5050_/A vssd1 vssd1 vccd1 vccd1 _5050_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4001_ _2896_/A _3935_/C _4288_/A vssd1 vssd1 vccd1 vccd1 _4001_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4606__A _5379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5952_ _6064_/CLK _5952_/D vssd1 vssd1 vccd1 vccd1 _5952_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_46_wb_clk_i_A clkbuf_3_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_18_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4903_ _5976_/Q _4859_/X _4869_/X _4902_/X vssd1 vssd1 vccd1 vccd1 _4903_/X sky130_fd_sc_hd__a211o_1
XFILLER_21_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5883_ _6027_/CLK _5883_/D vssd1 vssd1 vccd1 vccd1 _5883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4834_ _6087_/Q _4834_/B vssd1 vssd1 vccd1 vccd1 _4834_/X sky130_fd_sc_hd__or2_1
XFILLER_21_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3918__A1 _3037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4765_ _5401_/A _4602_/X _4756_/A vssd1 vssd1 vccd1 vccd1 _4765_/Y sky130_fd_sc_hd__a21oi_1
X_3716_ input6/X _5690_/Q _3735_/S vssd1 vssd1 vccd1 vccd1 _3716_/X sky130_fd_sc_hd__mux2_1
X_4696_ _5885_/Q _4653_/X _4694_/X _4695_/X vssd1 vssd1 vccd1 vccd1 _5885_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3647_ _5369_/A _5672_/Q _3651_/S vssd1 vssd1 vccd1 vccd1 _3648_/B sky130_fd_sc_hd__mux2_1
X_3578_ _5622_/A _5581_/A vssd1 vssd1 vccd1 vccd1 _5654_/B sky130_fd_sc_hd__nor2_1
XFILLER_88_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5317_ _5311_/Y _5312_/X _5316_/X _5266_/X vssd1 vssd1 vccd1 vccd1 _5317_/Y sky130_fd_sc_hd__o211ai_1
XANTENNA__5172__A _5638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5248_ _5248_/A _5248_/B vssd1 vssd1 vccd1 vccd1 _5269_/C sky130_fd_sc_hd__nor2_1
XFILLER_56_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5179_ _5056_/A _5990_/Q _5189_/S vssd1 vssd1 vccd1 vccd1 _5180_/B sky130_fd_sc_hd__mux2_1
XFILLER_56_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3420__A _5171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4251__A _4251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4334__B2 _6065_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4397__S _4397_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_435 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2880_ _2880_/A vssd1 vssd1 vccd1 vccd1 _3836_/A sky130_fd_sc_hd__buf_2
XFILLER_30_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4550_ _4550_/A _4550_/B vssd1 vssd1 vccd1 vccd1 _4550_/Y sky130_fd_sc_hd__nor2_1
X_4481_ _3553_/X _4530_/A _4480_/Y _5857_/Q vssd1 vssd1 vccd1 vccd1 _4481_/X sky130_fd_sc_hd__o31a_1
X_3501_ _3161_/A _3493_/X _3117_/Y _3500_/Y _3374_/A vssd1 vssd1 vccd1 vccd1 _3502_/B
+ sky130_fd_sc_hd__a32o_1
X_3432_ _4437_/B _3432_/B _2936_/A vssd1 vssd1 vccd1 vccd1 _3432_/X sky130_fd_sc_hd__or3b_1
XANTENNA__4325__A1 _3820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3363_ _3332_/X _3353_/X _3361_/X _3368_/C vssd1 vssd1 vccd1 vccd1 _3386_/A sky130_fd_sc_hd__o31a_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_41_wb_clk_i clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5983_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__3505__A _3668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5102_ _5102_/A vssd1 vssd1 vccd1 vccd1 _5535_/B sky130_fd_sc_hd__clkbuf_2
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3294_ _4217_/A vssd1 vssd1 vccd1 vccd1 _5241_/C sky130_fd_sc_hd__clkbuf_2
X_6082_ _6085_/CLK _6082_/D vssd1 vssd1 vccd1 vccd1 _6082_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5033_ _5942_/Q _5036_/C vssd1 vssd1 vccd1 vccd1 _5035_/A sky130_fd_sc_hd__and2_1
XFILLER_38_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_2_wb_clk_i_A clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_53_435 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5935_ _5959_/CLK _5935_/D vssd1 vssd1 vccd1 vccd1 _5935_/Q sky130_fd_sc_hd__dfxtp_1
X_5866_ _5874_/CLK _5866_/D vssd1 vssd1 vccd1 vccd1 _5866_/Q sky130_fd_sc_hd__dfxtp_1
X_4817_ _5897_/Q _4807_/X _4815_/X _4816_/X vssd1 vssd1 vccd1 vccd1 _5897_/D sky130_fd_sc_hd__a22o_1
X_5797_ _5959_/CLK _5797_/D vssd1 vssd1 vccd1 vccd1 _5797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4564__A1 _5874_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4748_ _5703_/Q _5680_/Q _4748_/S vssd1 vssd1 vccd1 vccd1 _4748_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4679_ _4779_/A vssd1 vssd1 vccd1 vccd1 _4719_/S sky130_fd_sc_hd__clkbuf_2
Xoutput59 _5886_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[73] sky130_fd_sc_hd__buf_2
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5987__D _5987_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3150__A _3391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_490 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3981_ _3994_/A _3981_/B vssd1 vssd1 vccd1 vccd1 _3982_/A sky130_fd_sc_hd__and2_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2932_ _6012_/Q _6011_/Q _6010_/Q vssd1 vssd1 vccd1 vccd1 _2942_/A sky130_fd_sc_hd__or3b_1
X_5720_ _5796_/CLK _5720_/D vssd1 vssd1 vccd1 vccd1 _5720_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4794__A1 _6059_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2863_ _2863_/A vssd1 vssd1 vccd1 vccd1 _2863_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5651_ _5389_/X _3576_/A _5650_/X _5172_/X vssd1 vssd1 vccd1 vccd1 _6136_/D sky130_fd_sc_hd__o211a_1
X_5582_ _5599_/B vssd1 vssd1 vccd1 vccd1 _5592_/B sky130_fd_sc_hd__clkbuf_1
X_4602_ _4716_/A vssd1 vssd1 vccd1 vccd1 _4602_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4533_ _4534_/B _4527_/X _4534_/A vssd1 vssd1 vccd1 vccd1 _4535_/A sky130_fd_sc_hd__a21oi_1
XFILLER_7_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_proj_example_181 vssd1 vssd1 vccd1 vccd1 user_proj_example_181/HI la_data_out[56]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_170 vssd1 vssd1 vccd1 vccd1 user_proj_example_170/HI la_data_out[45]
+ sky130_fd_sc_hd__conb_1
XFILLER_89_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4464_ _2944_/B _4464_/B vssd1 vssd1 vccd1 vccd1 _4464_/X sky130_fd_sc_hd__and2b_1
Xuser_proj_example_192 vssd1 vssd1 vccd1 vccd1 user_proj_example_192/HI la_data_out[99]
+ sky130_fd_sc_hd__conb_1
X_3415_ _3415_/A _3415_/B vssd1 vssd1 vccd1 vccd1 _3415_/Y sky130_fd_sc_hd__nand2_1
X_4395_ _4395_/A vssd1 vssd1 vccd1 vccd1 _5834_/D sky130_fd_sc_hd__clkbuf_1
X_3346_ _4235_/C _3346_/B _3518_/B vssd1 vssd1 vccd1 vccd1 _3346_/X sky130_fd_sc_hd__and3_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6134_ _6135_/CLK _6134_/D vssd1 vssd1 vccd1 vccd1 _6134_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6065_ _6067_/CLK _6065_/D vssd1 vssd1 vccd1 vccd1 _6065_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_85_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3277_ _4220_/A _3275_/X _3260_/X _3276_/Y _3161_/X vssd1 vssd1 vccd1 vccd1 _3277_/Y
+ sky130_fd_sc_hd__o221ai_1
X_5016_ _5937_/Q _5936_/Q _5853_/Q _5016_/D vssd1 vssd1 vccd1 vccd1 _5023_/C sky130_fd_sc_hd__and4_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5450__A _5581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4066__A _4203_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5918_ _5988_/CLK _5918_/D vssd1 vssd1 vccd1 vccd1 _5918_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4785__A1 _6058_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5431__C1 _5420_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5849_ _6131_/CLK _5849_/D vssd1 vssd1 vccd1 vccd1 _5849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5360__A input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input14_A la_data_in[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4776__A1 _6033_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5489__C1 _5488_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3200_ _6025_/Q _5944_/Q vssd1 vssd1 vccd1 vccd1 _3200_/Y sky130_fd_sc_hd__xnor2_1
X_4180_ _5796_/Q _4179_/X _4184_/S vssd1 vssd1 vccd1 vccd1 _4181_/A sky130_fd_sc_hd__mux2_1
X_3131_ _5870_/Q vssd1 vssd1 vccd1 vccd1 _4548_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_79_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3062_ _3389_/A vssd1 vssd1 vccd1 vccd1 _5297_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_67_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3964_ _3964_/A vssd1 vssd1 vccd1 vccd1 _3964_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4614__A _4883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2915_ _3322_/A _3439_/A _5228_/B vssd1 vssd1 vccd1 vccd1 _3448_/A sky130_fd_sc_hd__a21o_1
X_3895_ _6112_/Q _3894_/X _4041_/S vssd1 vssd1 vccd1 vccd1 _3895_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5703_ _5703_/CLK _5703_/D vssd1 vssd1 vccd1 vccd1 _5703_/Q sky130_fd_sc_hd__dfxtp_1
X_2846_ _5281_/A _3063_/C _2846_/C vssd1 vssd1 vccd1 vccd1 _3507_/A sky130_fd_sc_hd__nand3_1
X_5634_ _5360_/X _5623_/X _5633_/X _5627_/X vssd1 vssd1 vccd1 vccd1 _6116_/D sky130_fd_sc_hd__o211a_1
X_5565_ _5353_/X _5559_/X _5564_/X _5556_/X vssd1 vssd1 vccd1 vccd1 _6090_/D sky130_fd_sc_hd__o211a_1
X_4516_ _4516_/A vssd1 vssd1 vccd1 vccd1 _5862_/D sky130_fd_sc_hd__clkbuf_1
X_5496_ _6065_/Q _5505_/B vssd1 vssd1 vccd1 vccd1 _5496_/X sky130_fd_sc_hd__or2_1
X_4447_ _4447_/A _6123_/Q _4447_/C _4447_/D vssd1 vssd1 vccd1 vccd1 _4447_/X sky130_fd_sc_hd__or4_1
XANTENNA_input6_A la_data_in[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4378_ _5829_/Q _4376_/X _4391_/S vssd1 vssd1 vccd1 vccd1 _4379_/A sky130_fd_sc_hd__mux2_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6117_ _6117_/CLK _6117_/D vssd1 vssd1 vccd1 vccd1 _6117_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3329_ _3486_/A _3305_/X _3310_/X _3319_/X _3328_/X vssd1 vssd1 vccd1 vccd1 _3329_/Y
+ sky130_fd_sc_hd__o2111ai_2
XFILLER_58_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5180__A _5186_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6048_ _6048_/CLK _6048_/D vssd1 vssd1 vccd1 vccd1 _6048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5355__A _5391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4930__A1 _6036_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5249__B _5258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3680_ _3680_/A vssd1 vssd1 vccd1 vccd1 _5681_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_290 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2889__A _3873_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5350_ _5374_/B vssd1 vssd1 vccd1 vccd1 _5367_/B sky130_fd_sc_hd__clkbuf_1
X_5281_ _5281_/A _5281_/B vssd1 vssd1 vccd1 vccd1 _5281_/Y sky130_fd_sc_hd__nor2_1
X_4301_ _4233_/B _4294_/C _3260_/X vssd1 vssd1 vccd1 vccd1 _4307_/A sky130_fd_sc_hd__a21oi_1
X_4232_ _3346_/B _3518_/B _5257_/A vssd1 vssd1 vccd1 vccd1 _4233_/C sky130_fd_sc_hd__a21bo_1
XFILLER_4_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4163_ _5791_/Q _4162_/X _4167_/S vssd1 vssd1 vccd1 vccd1 _4164_/A sky130_fd_sc_hd__mux2_1
X_3114_ _3410_/A vssd1 vssd1 vccd1 vccd1 _3161_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_67_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4094_ _4094_/A vssd1 vssd1 vccd1 vccd1 _5771_/D sky130_fd_sc_hd__clkbuf_1
X_3045_ _3857_/B _3045_/B vssd1 vssd1 vccd1 vccd1 _3046_/B sky130_fd_sc_hd__nand2_1
XFILLER_82_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4996_ _4996_/A vssd1 vssd1 vccd1 vccd1 _5930_/D sky130_fd_sc_hd__clkbuf_1
X_3947_ _3966_/A _3947_/B vssd1 vssd1 vccd1 vccd1 _3948_/A sky130_fd_sc_hd__and2_1
X_3878_ _3896_/A _3875_/X _3877_/Y _4210_/A vssd1 vssd1 vccd1 vccd1 _3878_/X sky130_fd_sc_hd__a211o_1
X_2829_ _5872_/Q vssd1 vssd1 vccd1 vccd1 _5245_/A sky130_fd_sc_hd__clkbuf_2
X_5617_ _3611_/X _5602_/A _5616_/X _5612_/X vssd1 vssd1 vccd1 vccd1 _6110_/D sky130_fd_sc_hd__o211a_1
X_5548_ _3604_/X _5536_/X _5547_/X _5545_/X vssd1 vssd1 vccd1 vccd1 _6084_/D sky130_fd_sc_hd__o211a_1
X_5479_ _6059_/Q _5483_/B vssd1 vssd1 vccd1 vccd1 _5479_/X sky130_fd_sc_hd__or2_1
XFILLER_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xuser_proj_example_90 vssd1 vssd1 vccd1 vccd1 user_proj_example_90/HI io_oeb[8] sky130_fd_sc_hd__conb_1
XFILLER_86_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4903__A1 _5976_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4667__A0 _6119_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_36_wb_clk_i_A clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_60_341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4850_ _5955_/Q _4849_/X _4873_/S vssd1 vssd1 vccd1 vccd1 _4850_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3801_ _3161_/X _3493_/X _3260_/X _5846_/Q vssd1 vssd1 vccd1 vccd1 _3801_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5395__A1 _5393_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4781_ _4781_/A vssd1 vssd1 vccd1 vccd1 _4822_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_9_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3732_ _3732_/A _3732_/B vssd1 vssd1 vccd1 vccd1 _3733_/A sky130_fd_sc_hd__and2_1
X_3663_ _3666_/A _3663_/B vssd1 vssd1 vccd1 vccd1 _3664_/A sky130_fd_sc_hd__and2_1
X_5402_ _3582_/X _5387_/B _5401_/Y _5391_/X vssd1 vssd1 vccd1 vccd1 _6032_/D sky130_fd_sc_hd__o211a_1
X_5333_ _6066_/Q _6013_/Q _5336_/S vssd1 vssd1 vccd1 vccd1 _5333_/X sky130_fd_sc_hd__mux2_1
X_3594_ _5624_/A _5603_/A vssd1 vssd1 vccd1 vccd1 _3618_/B sky130_fd_sc_hd__nor2_1
XFILLER_87_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5264_ _5243_/A _5262_/X _5246_/A _3547_/A vssd1 vssd1 vccd1 vccd1 _5264_/X sky130_fd_sc_hd__a31o_1
X_4215_ _3880_/S _3432_/B _3851_/D _4214_/X vssd1 vssd1 vccd1 vccd1 _4215_/X sky130_fd_sc_hd__a31o_1
X_5195_ _5072_/A _5995_/Q _5198_/S vssd1 vssd1 vccd1 vccd1 _5196_/B sky130_fd_sc_hd__mux2_1
X_4146_ _5786_/Q _4145_/X _4150_/S vssd1 vssd1 vccd1 vccd1 _4147_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3881__A1 _5301_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4077_ _4077_/A vssd1 vssd1 vccd1 vccd1 _5766_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3028_ _4438_/A vssd1 vssd1 vccd1 vccd1 _4283_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_70_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4979_ _5925_/Q _4948_/X _4975_/X _5926_/Q vssd1 vssd1 vccd1 vccd1 _4979_/X sky130_fd_sc_hd__a31o_1
XFILLER_78_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3153__A _3375_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2992__A _3256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4000_ _5188_/A vssd1 vssd1 vccd1 vccd1 _4524_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5951_ _5959_/CLK _5951_/D vssd1 vssd1 vccd1 vccd1 _5951_/Q sky130_fd_sc_hd__dfxtp_1
X_4902_ _4870_/X _4900_/X _4901_/X _4875_/X vssd1 vssd1 vccd1 vccd1 _4902_/X sky130_fd_sc_hd__o211a_1
X_5882_ _6027_/CLK _5882_/D vssd1 vssd1 vccd1 vccd1 _5882_/Q sky130_fd_sc_hd__dfxtp_1
X_4833_ _6111_/Q _4831_/X _4873_/S vssd1 vssd1 vccd1 vccd1 _4833_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5368__A1 _5366_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4576__C1 _4460_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4764_ _6056_/Q _4757_/X _4716_/X _4763_/X vssd1 vssd1 vccd1 vccd1 _4764_/X sky130_fd_sc_hd__a211o_1
XANTENNA__4341__B _6041_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3715_ _3722_/S vssd1 vssd1 vccd1 vccd1 _3735_/S sky130_fd_sc_hd__clkbuf_2
X_4695_ _6025_/Q _4674_/X _4675_/X vssd1 vssd1 vccd1 vccd1 _4695_/X sky130_fd_sc_hd__o21a_1
XANTENNA__3238__A _6030_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3646_ _3646_/A vssd1 vssd1 vccd1 vccd1 _5671_/D sky130_fd_sc_hd__clkbuf_1
X_3577_ _3577_/A vssd1 vssd1 vccd1 vccd1 _5581_/A sky130_fd_sc_hd__clkbuf_2
X_5316_ _3491_/X _5257_/Y _5314_/Y _5315_/Y vssd1 vssd1 vccd1 vccd1 _5316_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5247_ _5247_/A _5247_/B vssd1 vssd1 vccd1 vccd1 _5258_/B sky130_fd_sc_hd__nor2_2
XFILLER_75_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5178_ _5178_/A vssd1 vssd1 vccd1 vccd1 _5989_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4129_ _5781_/Q _4128_/X _4133_/S vssd1 vssd1 vccd1 vccd1 _4130_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3606__A1 _3604_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5359__A1 _5357_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2987__A _3841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5363__A input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input44_A wbs_sel_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4707__A _4914_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5598__A1 _3563_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3500_ _3354_/X _3411_/B _3493_/A _3396_/Y vssd1 vssd1 vccd1 vccd1 _3500_/Y sky130_fd_sc_hd__o31ai_1
X_4480_ _4480_/A _4568_/B vssd1 vssd1 vccd1 vccd1 _4480_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__2897__A _5279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3431_ _3427_/X _3428_/X _3430_/X _3448_/A vssd1 vssd1 vccd1 vccd1 _3431_/X sky130_fd_sc_hd__a31o_1
XANTENNA__4588__S _4914_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3362_ _4206_/A _5243_/B vssd1 vssd1 vccd1 vccd1 _3368_/C sky130_fd_sc_hd__nor2_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5101_ _5075_/X _5080_/A _5100_/X _5098_/X vssd1 vssd1 vccd1 vccd1 _5962_/D sky130_fd_sc_hd__o211a_1
X_3293_ _3293_/A _4259_/B vssd1 vssd1 vccd1 vccd1 _3300_/B sky130_fd_sc_hd__nor2_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6081_ _6085_/CLK _6081_/D vssd1 vssd1 vccd1 vccd1 _6081_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_528 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5032_ _5036_/C _5032_/B vssd1 vssd1 vccd1 vccd1 _5941_/D sky130_fd_sc_hd__nor2_1
XANTENNA__5589__A1 _5386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4261__A1 _3880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5934_ _5959_/CLK _5934_/D vssd1 vssd1 vccd1 vccd1 _5934_/Q sky130_fd_sc_hd__dfxtp_1
X_5865_ _5874_/CLK _5865_/D vssd1 vssd1 vccd1 vccd1 _5865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5448__A _5579_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4816_ _6037_/Q _4803_/X _4804_/X vssd1 vssd1 vccd1 vccd1 _4816_/X sky130_fd_sc_hd__o21a_1
XFILLER_33_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4013__A1 _6089_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5796_ _5796_/CLK _5796_/D vssd1 vssd1 vccd1 vccd1 _5796_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5210__A0 _5059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4747_ _5890_/Q _4705_/X _4743_/X _4746_/X vssd1 vssd1 vccd1 vccd1 _5890_/D sky130_fd_sc_hd__a22o_1
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4678_ _5696_/Q _5673_/Q _4697_/S vssd1 vssd1 vccd1 vccd1 _4678_/X sky130_fd_sc_hd__mux2_1
X_3629_ _3632_/A _3629_/B vssd1 vssd1 vccd1 vccd1 _3630_/A sky130_fd_sc_hd__and2_1
Xoutput49 _5874_/Q vssd1 vssd1 vccd1 vccd1 io_out[0] sky130_fd_sc_hd__buf_2
XANTENNA__5183__A _5186_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5358__A _6019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5504__A1 _5360_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5093__A _5959_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3980_ _5731_/Q _3964_/X _3953_/A _5730_/Q vssd1 vssd1 vccd1 vccd1 _3981_/B sky130_fd_sc_hd__a22o_1
XFILLER_62_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2931_ _3429_/B _2931_/B vssd1 vssd1 vccd1 vccd1 _3047_/A sky130_fd_sc_hd__or2_1
XANTENNA__4794__A2 _4757_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5650_ _6136_/Q _5654_/B vssd1 vssd1 vccd1 vccd1 _5650_/X sky130_fd_sc_hd__or2_1
XFILLER_87_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2862_ _2941_/A _2931_/B vssd1 vssd1 vccd1 vccd1 _2863_/A sky130_fd_sc_hd__or2_1
X_4601_ _4869_/A vssd1 vssd1 vccd1 vccd1 _4716_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5581_ _5581_/A _5601_/B vssd1 vssd1 vccd1 vccd1 _5599_/B sky130_fd_sc_hd__nor2_1
X_4532_ _4534_/B _4527_/X _4536_/B _4531_/Y vssd1 vssd1 vccd1 vccd1 _5865_/D sky130_fd_sc_hd__o211a_1
X_4463_ _4463_/A vssd1 vssd1 vccd1 vccd1 _5850_/D sky130_fd_sc_hd__clkbuf_1
Xuser_proj_example_171 vssd1 vssd1 vccd1 vccd1 user_proj_example_171/HI la_data_out[46]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_160 vssd1 vssd1 vccd1 vccd1 user_proj_example_160/HI la_data_out[35]
+ sky130_fd_sc_hd__conb_1
X_3414_ _3075_/B _3410_/X _3413_/X vssd1 vssd1 vccd1 vccd1 _3415_/B sky130_fd_sc_hd__a21o_1
XANTENNA__4111__S _4116_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xuser_proj_example_182 vssd1 vssd1 vccd1 vccd1 user_proj_example_182/HI la_data_out[57]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_193 vssd1 vssd1 vccd1 vccd1 user_proj_example_193/HI la_data_out[100]
+ sky130_fd_sc_hd__conb_1
X_4394_ _5834_/Q _4393_/X _4397_/S vssd1 vssd1 vccd1 vccd1 _4395_/A sky130_fd_sc_hd__mux2_1
X_3345_ _3841_/A _5715_/Q vssd1 vssd1 vccd1 vccd1 _3518_/B sky130_fd_sc_hd__or2_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6133_ _6135_/CLK _6133_/D vssd1 vssd1 vccd1 vccd1 _6133_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3276_ _5818_/Q _3898_/A vssd1 vssd1 vccd1 vccd1 _3276_/Y sky130_fd_sc_hd__nor2_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6064_ _6064_/CLK _6064_/D vssd1 vssd1 vccd1 vccd1 _6064_/Q sky130_fd_sc_hd__dfxtp_1
X_5015_ _5015_/A vssd1 vssd1 vccd1 vccd1 _5936_/D sky130_fd_sc_hd__clkbuf_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5450__B _5471_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5917_ _5920_/CLK _5917_/D vssd1 vssd1 vccd1 vccd1 _5917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4785__A2 _4757_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5848_ _6122_/CLK _5848_/D vssd1 vssd1 vccd1 vccd1 _5848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5779_ _6117_/CLK _5779_/D vssd1 vssd1 vccd1 vccd1 _5779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_70 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5535__B _5535_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5254__C _5254_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3503__A3 _3891_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3130_ _5742_/Q vssd1 vssd1 vccd1 vccd1 _4562_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_67_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3061_ _3061_/A _3061_/B vssd1 vssd1 vccd1 vccd1 _3127_/B sky130_fd_sc_hd__or2_1
XANTENNA__3071__A _3071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3963_ _3979_/A _3963_/B vssd1 vssd1 vccd1 vccd1 _5726_/D sky130_fd_sc_hd__nor2_1
XFILLER_35_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2914_ _3312_/D _2949_/C _5816_/Q vssd1 vssd1 vccd1 vccd1 _5228_/B sky130_fd_sc_hd__nor3b_2
X_3894_ _3880_/S _3891_/Y _3892_/X _3893_/X _5768_/Q vssd1 vssd1 vccd1 vccd1 _3894_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_50_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5702_ _5702_/CLK _5702_/D vssd1 vssd1 vccd1 vccd1 _5702_/Q sky130_fd_sc_hd__dfxtp_1
X_2845_ _3389_/A _3373_/B vssd1 vssd1 vccd1 vccd1 _2846_/C sky130_fd_sc_hd__and2_1
X_5633_ _6116_/Q _5635_/B vssd1 vssd1 vccd1 vccd1 _5633_/X sky130_fd_sc_hd__or2_1
X_5564_ _6090_/Q _5570_/B vssd1 vssd1 vccd1 vccd1 _5564_/X sky130_fd_sc_hd__or2_1
X_4515_ _4970_/A _4515_/B _4515_/C vssd1 vssd1 vccd1 vccd1 _4516_/A sky130_fd_sc_hd__and3_1
X_5495_ _5511_/B vssd1 vssd1 vccd1 vccd1 _5505_/B sky130_fd_sc_hd__clkbuf_1
X_4446_ _3415_/A _3092_/C _4278_/X _4445_/Y _4466_/A vssd1 vssd1 vccd1 vccd1 _4446_/X
+ sky130_fd_sc_hd__a2111o_1
X_4377_ _4397_/S vssd1 vssd1 vccd1 vccd1 _4391_/S sky130_fd_sc_hd__clkbuf_2
X_3328_ _3483_/A _3328_/B _3327_/X vssd1 vssd1 vccd1 vccd1 _3328_/X sky130_fd_sc_hd__or3b_1
XANTENNA__5461__A _5461_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6116_ _6117_/CLK _6116_/D vssd1 vssd1 vccd1 vccd1 _6116_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3259_ _3466_/D vssd1 vssd1 vccd1 vccd1 _4322_/B sky130_fd_sc_hd__clkbuf_2
X_6047_ _6048_/CLK _6047_/D vssd1 vssd1 vccd1 vccd1 _6047_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5371__A _5391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_26_wb_clk_i_A clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_60_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4921__A2 _4623_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5280_ _5280_/A vssd1 vssd1 vccd1 vccd1 _5281_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4300_ _4315_/A _4300_/B vssd1 vssd1 vccd1 vccd1 _5810_/D sky130_fd_sc_hd__nor2_1
X_4231_ _4231_/A _4231_/B vssd1 vssd1 vccd1 vccd1 _4233_/B sky130_fd_sc_hd__nand2_1
XFILLER_67_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4162_ _5659_/Q _5790_/Q _4162_/S vssd1 vssd1 vccd1 vccd1 _4162_/X sky130_fd_sc_hd__mux2_1
X_3113_ _3508_/B _3507_/A vssd1 vssd1 vccd1 vccd1 _5287_/A sky130_fd_sc_hd__and2_1
XFILLER_67_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4093_ _5771_/Q _4092_/X _4097_/S vssd1 vssd1 vccd1 vccd1 _4094_/A sky130_fd_sc_hd__mux2_1
X_3044_ _3465_/C _2959_/C _3465_/B _3044_/D vssd1 vssd1 vccd1 vccd1 _3857_/B sky130_fd_sc_hd__and4bb_2
XFILLER_67_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4995_ _5000_/C _4995_/B _4995_/C vssd1 vssd1 vccd1 vccd1 _4996_/A sky130_fd_sc_hd__and3b_1
X_3946_ _5723_/Q _3932_/A _3945_/X _5722_/Q vssd1 vssd1 vccd1 vccd1 _3947_/B sky130_fd_sc_hd__a22o_1
X_3877_ _3017_/B _3876_/Y _3896_/A vssd1 vssd1 vccd1 vccd1 _3877_/Y sky130_fd_sc_hd__a21oi_1
X_2828_ hold1/A vssd1 vssd1 vccd1 vccd1 _3929_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__4360__A _4397_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5616_ _6110_/Q _5620_/B vssd1 vssd1 vccd1 vccd1 _5616_/X sky130_fd_sc_hd__or2_1
X_5547_ _6084_/Q _5549_/B vssd1 vssd1 vccd1 vccd1 _5547_/X sky130_fd_sc_hd__or2_1
XANTENNA__4912__A2 _5379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5478_ _3598_/X _5470_/X _5475_/X _5477_/X vssd1 vssd1 vccd1 vccd1 _6058_/D sky130_fd_sc_hd__o211a_1
X_4429_ _5974_/Q _5844_/Q _4432_/S vssd1 vssd1 vccd1 vccd1 _4429_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4676__A1 _6023_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_proj_example_91 vssd1 vssd1 vccd1 vccd1 user_proj_example_91/HI io_oeb[9] sky130_fd_sc_hd__conb_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5366__A _5366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5313__C1 _5258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_122 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3800_ _3800_/A _3800_/B vssd1 vssd1 vccd1 vccd1 _3800_/Y sky130_fd_sc_hd__nand2_1
X_4780_ _5659_/Q _4778_/X _4821_/S vssd1 vssd1 vccd1 vccd1 _4780_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3731_ _5369_/A _5695_/Q _3735_/S vssd1 vssd1 vccd1 vccd1 _3732_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_35_wb_clk_i clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6040_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_9_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3662_ _5386_/A _5676_/Q _3669_/S vssd1 vssd1 vccd1 vccd1 _3663_/B sky130_fd_sc_hd__mux2_1
X_5401_ _5401_/A _5401_/B vssd1 vssd1 vccd1 vccd1 _5401_/Y sky130_fd_sc_hd__nand2_1
X_3593_ _3593_/A vssd1 vssd1 vccd1 vccd1 _5603_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5332_ _6065_/Q _3423_/A _5337_/S _5331_/X vssd1 vssd1 vccd1 vccd1 _6013_/D sky130_fd_sc_hd__a31o_1
X_5263_ _5287_/C _5251_/X _5262_/X vssd1 vssd1 vccd1 vccd1 _5263_/X sky130_fd_sc_hd__o21a_1
XFILLER_87_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4214_ _3282_/A _3821_/A _3849_/C _3296_/B _3814_/B vssd1 vssd1 vccd1 vccd1 _4214_/X
+ sky130_fd_sc_hd__a32o_1
X_5194_ _5194_/A vssd1 vssd1 vccd1 vccd1 _5994_/D sky130_fd_sc_hd__clkbuf_1
X_4145_ _6136_/Q _5785_/Q _4145_/S vssd1 vssd1 vccd1 vccd1 _4145_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_423 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4076_ _5766_/Q _4075_/X _4080_/S vssd1 vssd1 vccd1 vccd1 _4077_/A sky130_fd_sc_hd__mux2_1
XFILLER_70_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3027_ _5871_/Q vssd1 vssd1 vccd1 vccd1 _4438_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3897__C _4259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4978_ _4972_/B _4976_/Y _4977_/X _4940_/X vssd1 vssd1 vccd1 vccd1 _5925_/D sky130_fd_sc_hd__o211a_1
XFILLER_51_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3929_ _3927_/Y _3929_/B _3929_/C vssd1 vssd1 vccd1 vccd1 _3939_/A sky130_fd_sc_hd__and3b_1
XANTENNA__5186__A _5186_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2992__B _3296_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_66 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3609__A _5295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4337__A0 _6068_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5534__C1 _5529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5950_ _5959_/CLK _5950_/D vssd1 vssd1 vccd1 vccd1 _5950_/Q sky130_fd_sc_hd__dfxtp_1
X_4901_ _5968_/Q _4917_/B vssd1 vssd1 vccd1 vccd1 _4901_/X sky130_fd_sc_hd__or2_1
X_5881_ _6024_/CLK _5881_/D vssd1 vssd1 vccd1 vccd1 _5881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4832_ _4883_/A vssd1 vssd1 vccd1 vccd1 _4873_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__3918__A3 _4322_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4763_ _4717_/X _4761_/X _4762_/X _4722_/X vssd1 vssd1 vccd1 vccd1 _4763_/X sky130_fd_sc_hd__o211a_1
X_3714_ _5343_/B _5201_/A vssd1 vssd1 vccd1 vccd1 _3722_/S sky130_fd_sc_hd__nand2_2
X_4694_ _6049_/Q _4654_/X _4664_/X _4693_/X vssd1 vssd1 vccd1 vccd1 _4694_/X sky130_fd_sc_hd__a211o_1
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3645_ _3648_/A _3645_/B vssd1 vssd1 vccd1 vccd1 _3646_/A sky130_fd_sc_hd__and2_1
X_3576_ _3576_/A vssd1 vssd1 vccd1 vccd1 _3576_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5315_ _5315_/A _5315_/B vssd1 vssd1 vccd1 vccd1 _5315_/Y sky130_fd_sc_hd__xnor2_1
X_5246_ _5246_/A _5246_/B vssd1 vssd1 vccd1 vccd1 _5251_/B sky130_fd_sc_hd__nor2_1
XANTENNA__3254__A _4251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5177_ _5186_/A _5177_/B vssd1 vssd1 vccd1 vccd1 _5178_/A sky130_fd_sc_hd__and2_1
XFILLER_28_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4128_ _6118_/Q _5780_/Q _4128_/S vssd1 vssd1 vccd1 vccd1 _4128_/X sky130_fd_sc_hd__mux2_1
X_4059_ _5761_/Q _4058_/X _4063_/S vssd1 vssd1 vccd1 vccd1 _4060_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_331 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input37_A la_data_in[61] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3430_ _3430_/A _3483_/B _3429_/X vssd1 vssd1 vccd1 vccd1 _3430_/X sky130_fd_sc_hd__or3b_1
X_3361_ _3291_/B _3356_/X _3520_/B _3360_/X vssd1 vssd1 vccd1 vccd1 _3361_/X sky130_fd_sc_hd__a211o_1
XANTENNA__3505__C _3505_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3074__A _3873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6080_ _6080_/CLK _6080_/D vssd1 vssd1 vccd1 vccd1 _6080_/Q sky130_fd_sc_hd__dfxtp_1
X_5100_ _5962_/Q _5100_/B vssd1 vssd1 vccd1 vccd1 _5100_/X sky130_fd_sc_hd__or2_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3292_ _3849_/A _3264_/A _3017_/B vssd1 vssd1 vccd1 vccd1 _4259_/B sky130_fd_sc_hd__o21ai_2
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5031_ _5941_/Q _5029_/A _5020_/X vssd1 vssd1 vccd1 vccd1 _5032_/B sky130_fd_sc_hd__o21ai_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3802__A _5976_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_50_wb_clk_i clkbuf_3_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6108_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_5933_ _5959_/CLK _5933_/D vssd1 vssd1 vccd1 vccd1 _5933_/Q sky130_fd_sc_hd__dfxtp_1
X_5864_ _5926_/CLK _5864_/D vssd1 vssd1 vccd1 vccd1 _5864_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5448__B _5469_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4815_ _6061_/Q _4808_/X _4767_/X _4814_/X vssd1 vssd1 vccd1 vccd1 _4815_/X sky130_fd_sc_hd__a211o_1
XANTENNA__3249__A _4436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4013__A2 _3061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5795_ _6112_/CLK _5795_/D vssd1 vssd1 vccd1 vccd1 _5795_/Q sky130_fd_sc_hd__dfxtp_1
X_4746_ _6030_/Q _4744_/X _4745_/X vssd1 vssd1 vccd1 vccd1 _4746_/X sky130_fd_sc_hd__o21a_1
X_4677_ _5883_/Q _4653_/X _4672_/X _4676_/X vssd1 vssd1 vccd1 vccd1 _5883_/D sky130_fd_sc_hd__a22o_1
X_3628_ input5/X _5666_/Q _3641_/S vssd1 vssd1 vccd1 vccd1 _3629_/B sky130_fd_sc_hd__mux2_1
X_3559_ _3546_/A _3547_/Y _3556_/B _3558_/X vssd1 vssd1 vccd1 vccd1 _5743_/D sky130_fd_sc_hd__a31o_1
XFILLER_0_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_367 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5229_ _5229_/A _5229_/B vssd1 vssd1 vccd1 vccd1 _5229_/Y sky130_fd_sc_hd__nor2_1
XFILLER_48_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4808__A _4859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4252__A2 _3842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3159__A _3873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2998__A _3481_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5374__A _6024_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5440__A1 _5363_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2930_ _3874_/A vssd1 vssd1 vccd1 vccd1 _3466_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_50_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2861_ _6012_/Q _6010_/Q _6011_/Q vssd1 vssd1 vccd1 vccd1 _2931_/B sky130_fd_sc_hd__or3b_1
XFILLER_62_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4600_ _4604_/A _4604_/B vssd1 vssd1 vccd1 vccd1 _4869_/A sky130_fd_sc_hd__nor2_2
X_5580_ _5580_/A vssd1 vssd1 vccd1 vccd1 _5580_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4531_ _4534_/B _4527_/X _4436_/A vssd1 vssd1 vccd1 vccd1 _4531_/Y sky130_fd_sc_hd__a21oi_1
X_4462_ _5847_/Q _5850_/Q _4462_/S vssd1 vssd1 vccd1 vccd1 _4463_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5284__A _5284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xuser_proj_example_172 vssd1 vssd1 vccd1 vccd1 user_proj_example_172/HI la_data_out[47]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_150 vssd1 vssd1 vccd1 vccd1 user_proj_example_150/HI la_data_out[25]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_161 vssd1 vssd1 vccd1 vccd1 user_proj_example_161/HI la_data_out[36]
+ sky130_fd_sc_hd__conb_1
XANTENNA__3506__A1 _3255_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3413_ _3391_/A _3522_/B _3274_/C _3349_/C _3412_/X vssd1 vssd1 vccd1 vccd1 _3413_/X
+ sky130_fd_sc_hd__a41o_1
Xuser_proj_example_183 vssd1 vssd1 vccd1 vccd1 user_proj_example_183/HI la_data_out[58]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_194 vssd1 vssd1 vccd1 vccd1 user_proj_example_194/HI la_data_out[101]
+ sky130_fd_sc_hd__conb_1
XANTENNA__4703__B1 _4623_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4393_ _6056_/Q _5833_/Q _4396_/S vssd1 vssd1 vccd1 vccd1 _4393_/X sky130_fd_sc_hd__mux2_1
X_6132_ _6132_/CLK _6132_/D vssd1 vssd1 vccd1 vccd1 _6132_/Q sky130_fd_sc_hd__dfxtp_1
X_3344_ _3853_/A _5715_/Q vssd1 vssd1 vccd1 vccd1 _3346_/B sky130_fd_sc_hd__nand2_1
XFILLER_58_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3275_ _5818_/Q vssd1 vssd1 vccd1 vccd1 _3275_/X sky130_fd_sc_hd__clkbuf_2
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6063_ _6064_/CLK _6063_/D vssd1 vssd1 vccd1 vccd1 _6063_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5014_ _5025_/B _5014_/B _5014_/C vssd1 vssd1 vccd1 vccd1 _5015_/A sky130_fd_sc_hd__and3_1
XANTENNA__3809__A2 _3497_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5431__A1 _5342_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5916_ _5920_/CLK _5916_/D vssd1 vssd1 vccd1 vccd1 _5916_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_407 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5847_ _6131_/CLK _5847_/D vssd1 vssd1 vccd1 vccd1 _5847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5778_ _6117_/CLK _5778_/D vssd1 vssd1 vccd1 vccd1 _5778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4729_ _6137_/Q _4727_/X _4770_/S vssd1 vssd1 vccd1 vccd1 _4729_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_307 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_16_wb_clk_i_A _5836_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5369__A _5369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3336__B _3481_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5489__A1 _3614_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_55_wb_clk_i_A clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_4_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output68_A _5895_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3060_ _2863_/X _2900_/Y _4210_/B _3059_/X _3272_/B vssd1 vssd1 vccd1 vccd1 _3061_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_63_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5279__A _5279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3962_ _5726_/Q _3932_/X _3961_/X vssd1 vssd1 vccd1 vccd1 _3963_/B sky130_fd_sc_hd__a21oi_1
X_5701_ _5702_/CLK _5701_/D vssd1 vssd1 vccd1 vccd1 _5701_/Q sky130_fd_sc_hd__dfxtp_1
X_3893_ _4437_/B _3878_/X _3867_/A _3111_/X vssd1 vssd1 vccd1 vccd1 _3893_/X sky130_fd_sc_hd__a211o_1
X_2913_ _5815_/Q vssd1 vssd1 vccd1 vccd1 _3312_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_2844_ _6006_/Q _6007_/Q vssd1 vssd1 vccd1 vccd1 _3373_/B sky130_fd_sc_hd__and2b_1
X_5632_ _5357_/X _5623_/X _5631_/X _5627_/X vssd1 vssd1 vccd1 vccd1 _6115_/D sky130_fd_sc_hd__o211a_1
X_5563_ _5342_/X _5559_/X _5562_/X _5556_/X vssd1 vssd1 vccd1 vccd1 _6089_/D sky130_fd_sc_hd__o211a_1
X_4514_ _5862_/Q _4514_/B vssd1 vssd1 vccd1 vccd1 _4515_/C sky130_fd_sc_hd__nand2_1
X_5494_ _5537_/B _5624_/B vssd1 vssd1 vccd1 vccd1 _5511_/B sky130_fd_sc_hd__nor2_1
X_4445_ _3802_/B _3493_/A _4444_/X vssd1 vssd1 vccd1 vccd1 _4445_/Y sky130_fd_sc_hd__o21ai_1
X_4376_ _6051_/Q _5828_/Q _4380_/S vssd1 vssd1 vccd1 vccd1 _4376_/X sky130_fd_sc_hd__mux2_1
XFILLER_85_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3327_ _2997_/A _3159_/B _4438_/A vssd1 vssd1 vccd1 vccd1 _3327_/X sky130_fd_sc_hd__mux2_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6115_ _6115_/CLK _6115_/D vssd1 vssd1 vccd1 vccd1 _6115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3258_ _3851_/C vssd1 vssd1 vccd1 vccd1 _3466_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_58_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6046_ _6048_/CLK _6046_/D vssd1 vssd1 vccd1 vccd1 _6046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3189_ _5923_/Q _5914_/Q vssd1 vssd1 vccd1 vccd1 _3189_/Y sky130_fd_sc_hd__nand2_1
XFILLER_54_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4915__A0 _5954_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2979__C _4220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5643__A1 _5373_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4230_ _5327_/B _3316_/X _3318_/X _4229_/Y vssd1 vssd1 vccd1 vccd1 _4231_/B sky130_fd_sc_hd__a31o_1
XFILLER_4_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5562__A _6089_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4161_ _4161_/A vssd1 vssd1 vccd1 vccd1 _5790_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3082__A _3480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3112_ _3820_/A _3111_/X _3476_/C _3283_/B vssd1 vssd1 vccd1 vccd1 _3112_/X sky130_fd_sc_hd__a31o_1
X_4092_ _5957_/Q _5770_/Q _4092_/S vssd1 vssd1 vccd1 vccd1 _4092_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5634__A1 _5360_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3043_ _3035_/X _3037_/Y _3042_/X vssd1 vssd1 vccd1 vccd1 _3043_/X sky130_fd_sc_hd__o21a_1
XFILLER_48_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4994_ _5929_/Q _4993_/C _5930_/Q vssd1 vssd1 vccd1 vccd1 _4995_/C sky130_fd_sc_hd__a21o_1
X_3945_ _3952_/A vssd1 vssd1 vccd1 vccd1 _3945_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3876_ _3849_/A _3264_/A _3845_/C vssd1 vssd1 vccd1 vccd1 _3876_/Y sky130_fd_sc_hd__o21ai_1
X_5615_ _3607_/X _5602_/X _5614_/X _5612_/X vssd1 vssd1 vccd1 vccd1 _6109_/D sky130_fd_sc_hd__o211a_1
X_5546_ _3601_/X _5536_/X _5543_/X _5545_/X vssd1 vssd1 vccd1 vccd1 _6083_/D sky130_fd_sc_hd__o211a_1
X_5477_ _5529_/A vssd1 vssd1 vccd1 vccd1 _5477_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3581__C1 _3221_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4428_ _4428_/A vssd1 vssd1 vccd1 vccd1 _5844_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3884__A0 _6104_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4359_ _6046_/Q _5823_/Q _4363_/S vssd1 vssd1 vccd1 vccd1 _4359_/X sky130_fd_sc_hd__mux2_1
Xuser_proj_example_92 vssd1 vssd1 vccd1 vccd1 user_proj_example_92/HI io_oeb[10] sky130_fd_sc_hd__conb_1
XFILLER_58_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6029_ _6031_/CLK _6029_/D vssd1 vssd1 vccd1 vccd1 _6029_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_5_wb_clk_i clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6091_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_73_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3720__A _5875_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4052__A0 _6101_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3730_ _3730_/A vssd1 vssd1 vccd1 vccd1 _5694_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3661_ _3661_/A vssd1 vssd1 vccd1 vccd1 _5675_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5400_ _3563_/X _5387_/B _5399_/X _5391_/X vssd1 vssd1 vccd1 vccd1 _6031_/D sky130_fd_sc_hd__o211a_1
X_3592_ _3592_/A vssd1 vssd1 vccd1 vccd1 _3592_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5331_ _5337_/S _6013_/Q vssd1 vssd1 vccd1 vccd1 _5331_/X sky130_fd_sc_hd__and2b_1
X_5262_ _5294_/S vssd1 vssd1 vccd1 vccd1 _5262_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4213_ _3037_/A _3042_/X _3839_/D _4212_/X vssd1 vssd1 vccd1 vccd1 _4213_/X sky130_fd_sc_hd__a31o_1
XFILLER_68_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5193_ _5204_/A _5193_/B vssd1 vssd1 vccd1 vccd1 _5194_/A sky130_fd_sc_hd__and2_1
XFILLER_68_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4144_ _4144_/A vssd1 vssd1 vccd1 vccd1 _5785_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_435 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4075_ _6109_/Q _5765_/Q _4075_/S vssd1 vssd1 vccd1 vccd1 _4075_/X sky130_fd_sc_hd__mux2_1
X_3026_ _3482_/A vssd1 vssd1 vccd1 vccd1 _3897_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__3897__D _3897_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4977_ _4948_/X _4975_/X _5925_/Q vssd1 vssd1 vccd1 vccd1 _4977_/X sky130_fd_sc_hd__a21o_1
X_3928_ _3928_/A _3928_/B _3335_/C vssd1 vssd1 vccd1 vccd1 _3929_/C sky130_fd_sc_hd__or3b_1
X_3859_ _4280_/A _6005_/Q _3859_/C _3873_/D vssd1 vssd1 vccd1 vccd1 _3874_/B sky130_fd_sc_hd__or4_1
XFILLER_50_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5529_ _5529_/A vssd1 vssd1 vccd1 vccd1 _5529_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_59_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3715__A _3722_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_148 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5231__C1 _3331_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5377__A _5581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3625__A _3794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output50_A _5877_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4900_ _5960_/Q _4899_/X _4916_/S vssd1 vssd1 vccd1 vccd1 _4900_/X sky130_fd_sc_hd__mux2_1
X_5880_ _6024_/CLK _5880_/D vssd1 vssd1 vccd1 vccd1 _5880_/Q sky130_fd_sc_hd__dfxtp_1
X_4831_ _5664_/Q _4829_/X _4872_/S vssd1 vssd1 vccd1 vccd1 _4831_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4762_ _6080_/Q _4783_/B vssd1 vssd1 vccd1 vccd1 _4762_/X sky130_fd_sc_hd__or2_1
X_3713_ _3794_/A _3798_/C vssd1 vssd1 vccd1 vccd1 _5201_/A sky130_fd_sc_hd__and2_2
X_4693_ _4665_/X _4690_/X _4692_/X _4670_/X vssd1 vssd1 vccd1 vccd1 _4693_/X sky130_fd_sc_hd__o211a_1
X_3644_ _5366_/A _5671_/Q _3651_/S vssd1 vssd1 vccd1 vccd1 _3645_/B sky130_fd_sc_hd__mux2_1
X_3575_ _5622_/A _5579_/A vssd1 vssd1 vccd1 vccd1 _3576_/A sky130_fd_sc_hd__or2_1
X_5314_ _3486_/A _2863_/X _5313_/X _5301_/A vssd1 vssd1 vccd1 vccd1 _5314_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_0_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5245_ _5245_/A _5245_/B vssd1 vssd1 vccd1 vccd1 _5246_/B sky130_fd_sc_hd__nor2_1
X_5176_ _5045_/A _5989_/Q _5189_/S vssd1 vssd1 vccd1 vccd1 _5177_/B sky130_fd_sc_hd__mux2_1
XFILLER_28_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4366__A _4366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4127_ _4127_/A vssd1 vssd1 vccd1 vccd1 _5780_/D sky130_fd_sc_hd__clkbuf_1
X_4058_ _6103_/Q _5760_/Q _4058_/S vssd1 vssd1 vccd1 vccd1 _4058_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3009_ _3824_/A _5720_/Q vssd1 vssd1 vccd1 vccd1 _3017_/B sky130_fd_sc_hd__xnor2_2
XFILLER_61_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4276__A _4276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3360_ _3440_/A _3360_/B _3821_/C vssd1 vssd1 vccd1 vccd1 _3360_/X sky130_fd_sc_hd__and3_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3291_ _3440_/A _3291_/B _3291_/C vssd1 vssd1 vccd1 vccd1 _3291_/X sky130_fd_sc_hd__and3_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ _5941_/Q _5940_/Q _5030_/C vssd1 vssd1 vccd1 vccd1 _5036_/C sky130_fd_sc_hd__and3_1
XANTENNA__4494__B1 _3999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3090__A _3375_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3802__B _3802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5932_ _5959_/CLK _5932_/D vssd1 vssd1 vccd1 vccd1 _5932_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5863_ _5926_/CLK _5863_/D vssd1 vssd1 vccd1 vccd1 _5863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4814_ _4768_/X _4812_/X _4813_/X _4773_/X vssd1 vssd1 vccd1 vccd1 _4814_/X sky130_fd_sc_hd__o211a_1
XFILLER_21_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5794_ _6109_/CLK _5794_/D vssd1 vssd1 vccd1 vccd1 _5794_/Q sky130_fd_sc_hd__dfxtp_1
X_4745_ _4855_/A vssd1 vssd1 vccd1 vccd1 _4745_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4676_ _6023_/Q _4674_/X _4675_/X vssd1 vssd1 vccd1 vccd1 _4676_/X sky130_fd_sc_hd__o21a_1
XANTENNA__2980__B1 _3518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3265__A _3854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3627_ _3651_/S vssd1 vssd1 vccd1 vccd1 _3641_/S sky130_fd_sc_hd__clkbuf_2
X_3558_ _5744_/Q _4331_/B _3412_/X _5743_/Q vssd1 vssd1 vccd1 vccd1 _3558_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3524__A2 _2955_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3489_ _3489_/A _3489_/B _3488_/X vssd1 vssd1 vccd1 vccd1 _3489_/X sky130_fd_sc_hd__or3b_1
XFILLER_88_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5228_ _5234_/A _5228_/B _4466_/B vssd1 vssd1 vccd1 vccd1 _5229_/A sky130_fd_sc_hd__or3b_1
XFILLER_56_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5159_ _5059_/X _5149_/X _5156_/X _5158_/X vssd1 vssd1 vccd1 vccd1 _5981_/D sky130_fd_sc_hd__o211a_1
XFILLER_29_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4824__A _4824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3159__B _3159_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_45_wb_clk_i_A clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__5390__A _6028_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5425__C1 _5420_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2860_ _3389_/A _5277_/A _6007_/Q _5277_/C vssd1 vssd1 vccd1 vccd1 _2941_/A sky130_fd_sc_hd__nand4_2
X_4530_ _4530_/A _4538_/B _4527_/X vssd1 vssd1 vccd1 vccd1 _4536_/B sky130_fd_sc_hd__or3b_1
XFILLER_7_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4461_ _5269_/A _4456_/X _4457_/X _4460_/X vssd1 vssd1 vccd1 vccd1 _5849_/D sky130_fd_sc_hd__o211a_1
Xuser_proj_example_140 vssd1 vssd1 vccd1 vccd1 user_proj_example_140/HI la_data_out[15]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_151 vssd1 vssd1 vccd1 vccd1 user_proj_example_151/HI la_data_out[26]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_162 vssd1 vssd1 vccd1 vccd1 user_proj_example_162/HI la_data_out[37]
+ sky130_fd_sc_hd__conb_1
X_3412_ _3412_/A vssd1 vssd1 vccd1 vccd1 _3412_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__3506__A2 _4409_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xuser_proj_example_184 vssd1 vssd1 vccd1 vccd1 user_proj_example_184/HI la_data_out[59]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_173 vssd1 vssd1 vccd1 vccd1 user_proj_example_173/HI la_data_out[48]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_195 vssd1 vssd1 vccd1 vccd1 user_proj_example_195/HI la_data_out[102]
+ sky130_fd_sc_hd__conb_1
XANTENNA__4703__A1 _5384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6131_ _6131_/CLK _6131_/D vssd1 vssd1 vccd1 vccd1 _6131_/Q sky130_fd_sc_hd__dfxtp_1
X_4392_ _4392_/A vssd1 vssd1 vccd1 vccd1 _5833_/D sky130_fd_sc_hd__clkbuf_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3343_ _6126_/Q vssd1 vssd1 vccd1 vccd1 _4235_/C sky130_fd_sc_hd__clkbuf_2
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3274_ _3820_/A _3274_/B _3274_/C _3423_/C vssd1 vssd1 vccd1 vccd1 _3274_/X sky130_fd_sc_hd__or4b_1
XANTENNA__4467__B1 _5803_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6062_ _6088_/CLK _6062_/D vssd1 vssd1 vccd1 vccd1 _6062_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5013_ _4946_/C _4982_/C _5936_/Q vssd1 vssd1 vccd1 vccd1 _5014_/C sky130_fd_sc_hd__a21o_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5915_ _5920_/CLK _5915_/D vssd1 vssd1 vccd1 vccd1 _5915_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_419 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5846_ _5944_/CLK _5846_/D vssd1 vssd1 vccd1 vccd1 _5846_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2989_ _3389_/A _5277_/A _6007_/Q _3407_/A vssd1 vssd1 vccd1 vccd1 _2990_/B sky130_fd_sc_hd__or4_1
X_5777_ _5777_/CLK _5777_/D vssd1 vssd1 vccd1 vccd1 _5777_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5475__A _6058_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4728_ _4779_/A vssd1 vssd1 vccd1 vccd1 _4770_/S sky130_fd_sc_hd__clkbuf_2
X_4659_ _6070_/Q _4683_/B vssd1 vssd1 vccd1 vccd1 _4659_/X sky130_fd_sc_hd__or2_1
XFILLER_1_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4819__A _4870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5655__C1 _5172_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_319 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_1_wb_clk_i_A clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_4_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_29_wb_clk_i clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5944_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_35_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3961_ _5725_/Q _3941_/X _3953_/X _3960_/Y vssd1 vssd1 vccd1 vccd1 _3961_/X sky130_fd_sc_hd__o211a_1
X_2912_ _3288_/C vssd1 vssd1 vccd1 vccd1 _3439_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5700_ _5702_/CLK _5700_/D vssd1 vssd1 vccd1 vccd1 _5700_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3892_ _3410_/A _3287_/X _3466_/D _5768_/Q vssd1 vssd1 vccd1 vccd1 _3892_/X sky130_fd_sc_hd__a31o_1
X_2843_ _6009_/Q vssd1 vssd1 vccd1 vccd1 _3389_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5295__A _5295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5631_ _6115_/Q _5635_/B vssd1 vssd1 vccd1 vccd1 _5631_/X sky130_fd_sc_hd__or2_1
X_5562_ _6089_/Q _5570_/B vssd1 vssd1 vccd1 vccd1 _5562_/X sky130_fd_sc_hd__or2_1
X_4513_ _4518_/C _4518_/D _4504_/Y _5862_/Q vssd1 vssd1 vccd1 vccd1 _4515_/B sky130_fd_sc_hd__a31o_1
X_5493_ _5493_/A vssd1 vssd1 vccd1 vccd1 _5493_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4444_ _3423_/A _3081_/B _4321_/S _4239_/A vssd1 vssd1 vccd1 vccd1 _4444_/X sky130_fd_sc_hd__o22a_1
X_4375_ _4375_/A vssd1 vssd1 vccd1 vccd1 _5828_/D sky130_fd_sc_hd__clkbuf_1
X_3326_ _3326_/A _3430_/A vssd1 vssd1 vccd1 vccd1 _3328_/B sky130_fd_sc_hd__nand2_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6114_ _6115_/CLK _6114_/D vssd1 vssd1 vccd1 vccd1 _6114_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6045_ _6048_/CLK _6045_/D vssd1 vssd1 vccd1 vccd1 _6045_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3112__B1 _3283_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3257_ _3257_/A vssd1 vssd1 vccd1 vccd1 _3851_/C sky130_fd_sc_hd__clkbuf_2
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_371 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3188_ _5924_/Q _4939_/A _4928_/A _5919_/Q vssd1 vssd1 vccd1 vccd1 _3188_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_54_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5829_ _6050_/CLK _5829_/D vssd1 vssd1 vccd1 vccd1 _5829_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3718__A _5171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_127 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input12_A la_data_in[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4459__A _5408_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4160_ _5790_/Q _4159_/X _4167_/S vssd1 vssd1 vccd1 vccd1 _4161_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3111_ _3821_/A vssd1 vssd1 vccd1 vccd1 _3111_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4091_ _4091_/A vssd1 vssd1 vccd1 vccd1 _5770_/D sky130_fd_sc_hd__clkbuf_1
X_3042_ _3042_/A vssd1 vssd1 vccd1 vccd1 _3042_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_500 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5398__A1 _5396_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4993_ _5930_/Q _5929_/Q _4993_/C vssd1 vssd1 vccd1 vccd1 _5000_/C sky130_fd_sc_hd__and3_1
X_3944_ _3954_/A _3940_/B vssd1 vssd1 vccd1 vccd1 _3952_/A sky130_fd_sc_hd__or2b_1
X_3875_ _3874_/A _3464_/Y _3872_/X _3874_/X vssd1 vssd1 vccd1 vccd1 _3875_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_31_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5614_ _6109_/Q _5614_/B vssd1 vssd1 vccd1 vccd1 _5614_/X sky130_fd_sc_hd__or2_1
X_5545_ _5597_/A vssd1 vssd1 vccd1 vccd1 _5545_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5476_ _5544_/A vssd1 vssd1 vccd1 vccd1 _5529_/A sky130_fd_sc_hd__buf_2
X_4427_ _5844_/Q _4426_/X _4433_/S vssd1 vssd1 vccd1 vccd1 _4428_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input4_A la_data_in[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4358_ _4358_/A vssd1 vssd1 vccd1 vccd1 _5823_/D sky130_fd_sc_hd__clkbuf_1
Xuser_proj_example_93 vssd1 vssd1 vccd1 vccd1 user_proj_example_93/HI io_oeb[11] sky130_fd_sc_hd__conb_1
XFILLER_86_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3309_ _5255_/A _3054_/A _3037_/B _3466_/A vssd1 vssd1 vccd1 vccd1 _3310_/B sky130_fd_sc_hd__o22a_1
X_4289_ _6130_/Q _3349_/C _3341_/B _3350_/A _4447_/A vssd1 vssd1 vccd1 vccd1 _4289_/Y
+ sky130_fd_sc_hd__a221oi_1
XFILLER_58_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6028_ _6031_/CLK _6028_/D vssd1 vssd1 vccd1 vccd1 _6028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4832__A _4883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5313__B2 _4259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3660_ _3666_/A _3660_/B vssd1 vssd1 vccd1 vccd1 _3661_/A sky130_fd_sc_hd__and2_1
XANTENNA__5552__A1 _3611_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3591_ _5622_/A _5601_/A vssd1 vssd1 vccd1 vccd1 _3592_/A sky130_fd_sc_hd__or2_1
X_5330_ _5327_/A _5266_/X _5329_/X vssd1 vssd1 vccd1 vccd1 _6012_/D sky130_fd_sc_hd__o21ba_1
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5261_ _5261_/A _5261_/B _5261_/C vssd1 vssd1 vccd1 vccd1 _5294_/S sky130_fd_sc_hd__nor3_2
X_4212_ _4287_/A _3839_/B _4210_/Y _4211_/X _3335_/X vssd1 vssd1 vccd1 vccd1 _4212_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_87_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_44_wb_clk_i clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6003_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_5192_ _5069_/A _5994_/Q _5198_/S vssd1 vssd1 vccd1 vccd1 _5193_/B sky130_fd_sc_hd__mux2_1
XFILLER_68_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4143_ _5785_/Q _4142_/X _4150_/S vssd1 vssd1 vccd1 vccd1 _4144_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4074_ _4074_/A vssd1 vssd1 vccd1 vccd1 _5765_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3025_ _3853_/A vssd1 vssd1 vccd1 vccd1 _3482_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4976_ _5925_/Q _4975_/X _4948_/X vssd1 vssd1 vccd1 vccd1 _4976_/Y sky130_fd_sc_hd__a21boi_1
X_3927_ _5256_/B _6121_/Q vssd1 vssd1 vccd1 vccd1 _3927_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3858_ _3858_/A _4471_/A _3042_/A _3839_/D vssd1 vssd1 vccd1 vccd1 _3861_/A sky130_fd_sc_hd__or4bb_1
X_3789_ _3966_/A _3789_/B vssd1 vssd1 vccd1 vccd1 _3790_/A sky130_fd_sc_hd__and2_1
X_5528_ _6078_/Q _5533_/B vssd1 vssd1 vccd1 vccd1 _5528_/X sky130_fd_sc_hd__or2_1
X_5459_ _5389_/X _5449_/X _5458_/X _5446_/X vssd1 vssd1 vccd1 vccd1 _6052_/D sky130_fd_sc_hd__o211a_1
XFILLER_1_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_480 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5377__B _5405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5534__A1 _3582_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3906__A _4210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3625__B _4645_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4830_ _4881_/A vssd1 vssd1 vccd1 vccd1 _4872_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_45_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4761_ _6104_/Q _4760_/X _4771_/S vssd1 vssd1 vccd1 vccd1 _4761_/X sky130_fd_sc_hd__mux2_1
X_3712_ _4594_/A _3712_/B _4594_/B vssd1 vssd1 vccd1 vccd1 _3798_/C sky130_fd_sc_hd__nor3_1
X_4692_ _6073_/Q _4732_/B vssd1 vssd1 vccd1 vccd1 _4692_/X sky130_fd_sc_hd__or2_1
XANTENNA__4328__A2 _4327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5525__A1 _5389_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3643_ _3643_/A vssd1 vssd1 vccd1 vccd1 _5670_/D sky130_fd_sc_hd__clkbuf_1
X_5313_ _3466_/C _3047_/X _3407_/A _4259_/A _5258_/B vssd1 vssd1 vccd1 vccd1 _5313_/X
+ sky130_fd_sc_hd__o221a_1
X_3574_ _3577_/A vssd1 vssd1 vccd1 vccd1 _5579_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_88_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5244_ _5244_/A _5244_/B _5271_/B vssd1 vssd1 vccd1 vccd1 _5246_/A sky130_fd_sc_hd__or3b_1
X_5175_ _5198_/S vssd1 vssd1 vccd1 vccd1 _5189_/S sky130_fd_sc_hd__clkbuf_2
X_4126_ _5780_/Q _4125_/X _4133_/S vssd1 vssd1 vccd1 vccd1 _4127_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4057_ _4057_/A vssd1 vssd1 vccd1 vccd1 _5760_/D sky130_fd_sc_hd__clkbuf_1
X_3008_ _3842_/A _3293_/A _3007_/X vssd1 vssd1 vccd1 vccd1 _3010_/B sky130_fd_sc_hd__o21ai_1
XFILLER_71_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_480 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5213__A0 _5062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4959_ _4966_/A _4959_/B vssd1 vssd1 vccd1 vccd1 _5920_/D sky130_fd_sc_hd__nor2_1
XFILLER_61_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3726__A _3732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_35_wb_clk_i_A clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_10_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3461__A _3854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_414 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_7__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3290_ _3482_/A _3287_/X _4470_/C _3849_/B _3897_/B vssd1 vssd1 vccd1 vccd1 _3291_/C
+ sky130_fd_sc_hd__a32o_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5931_ _5959_/CLK _5931_/D vssd1 vssd1 vccd1 vccd1 _5931_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5862_ _5926_/CLK _5862_/D vssd1 vssd1 vccd1 vccd1 _5862_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4406__S _4409_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4813_ _6085_/Q _4834_/B vssd1 vssd1 vccd1 vccd1 _4813_/X sky130_fd_sc_hd__or2_1
X_5793_ _6109_/CLK _5793_/D vssd1 vssd1 vccd1 vccd1 _5793_/Q sky130_fd_sc_hd__dfxtp_1
X_4744_ _5403_/B vssd1 vssd1 vccd1 vccd1 _4744_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4675_ _4855_/A vssd1 vssd1 vccd1 vccd1 _4675_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3626_ _5343_/B _5174_/A vssd1 vssd1 vccd1 vccd1 _3651_/S sky130_fd_sc_hd__nand2_2
X_3557_ _3553_/X _4530_/A _3556_/Y _3221_/X vssd1 vssd1 vccd1 vccd1 _5742_/D sky130_fd_sc_hd__o31a_1
X_3488_ _3468_/X _3479_/X _3487_/X _3269_/X vssd1 vssd1 vccd1 vccd1 _3488_/X sky130_fd_sc_hd__a31o_1
X_5227_ _5227_/A vssd1 vssd1 vccd1 vccd1 _6004_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4377__A _4397_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5158_ _5391_/A vssd1 vssd1 vccd1 vccd1 _5158_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4109_ _4109_/A vssd1 vssd1 vccd1 vccd1 _5775_/D sky130_fd_sc_hd__clkbuf_1
X_5089_ _5957_/Q _5093_/B vssd1 vssd1 vccd1 vccd1 _5089_/X sky130_fd_sc_hd__or2_1
XFILLER_72_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input42_A wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xuser_proj_example_130 vssd1 vssd1 vccd1 vccd1 user_proj_example_130/HI la_data_out[5]
+ sky130_fd_sc_hd__conb_1
X_4460_ _5067_/A vssd1 vssd1 vccd1 vccd1 _4460_/X sky130_fd_sc_hd__buf_2
Xuser_proj_example_141 vssd1 vssd1 vccd1 vccd1 user_proj_example_141/HI la_data_out[16]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_152 vssd1 vssd1 vccd1 vccd1 user_proj_example_152/HI la_data_out[27]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_163 vssd1 vssd1 vccd1 vccd1 user_proj_example_163/HI la_data_out[38]
+ sky130_fd_sc_hd__conb_1
X_3411_ _3929_/B _3411_/B vssd1 vssd1 vccd1 vccd1 _3412_/A sky130_fd_sc_hd__nor2_1
XFILLER_7_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_proj_example_185 vssd1 vssd1 vccd1 vccd1 user_proj_example_185/HI la_data_out[60]
+ sky130_fd_sc_hd__conb_1
X_4391_ _5833_/Q _4390_/X _4391_/S vssd1 vssd1 vccd1 vccd1 _4392_/A sky130_fd_sc_hd__mux2_1
Xuser_proj_example_174 vssd1 vssd1 vccd1 vccd1 user_proj_example_174/HI la_data_out[49]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_196 vssd1 vssd1 vccd1 vccd1 user_proj_example_196/HI la_data_out[103]
+ sky130_fd_sc_hd__conb_1
X_6130_ _6130_/CLK _6130_/D vssd1 vssd1 vccd1 vccd1 _6130_/Q sky130_fd_sc_hd__dfxtp_1
X_3342_ _6129_/Q _4239_/B vssd1 vssd1 vccd1 vccd1 _3342_/X sky130_fd_sc_hd__and2_1
XANTENNA__5581__A _5581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4909__B _4917_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3273_ _3081_/X _3082_/Y _5339_/S vssd1 vssd1 vccd1 vccd1 _4233_/A sky130_fd_sc_hd__o21ai_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6061_ _6088_/CLK _6061_/D vssd1 vssd1 vccd1 vccd1 _6061_/Q sky130_fd_sc_hd__dfxtp_1
X_5012_ _5012_/A _5012_/B _4972_/A vssd1 vssd1 vccd1 vccd1 _5014_/B sky130_fd_sc_hd__or3b_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_203 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5914_ _5914_/CLK _5914_/D vssd1 vssd1 vccd1 vccd1 _5914_/Q sky130_fd_sc_hd__dfxtp_1
X_5845_ _5944_/CLK _5845_/D vssd1 vssd1 vccd1 vccd1 _5845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2988_ _3518_/A _3116_/A vssd1 vssd1 vccd1 vccd1 _3350_/B sky130_fd_sc_hd__nor2_1
X_5776_ _5777_/CLK _5776_/D vssd1 vssd1 vccd1 vccd1 _5776_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4727_ _5701_/Q _5678_/Q _4748_/S vssd1 vssd1 vccd1 vccd1 _4727_/X sky130_fd_sc_hd__mux2_1
X_4658_ _6094_/Q _4657_/X _4668_/S vssd1 vssd1 vccd1 vccd1 _4658_/X sky130_fd_sc_hd__mux2_1
X_3609_ _5295_/A vssd1 vssd1 vccd1 vccd1 _3609_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__5352__C1 _5169_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4589_ _4881_/A vssd1 vssd1 vccd1 vccd1 _4779_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_1_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3723__B _5875_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4394__A0 _5834_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4918__C1 _5469_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4449__A1 _3820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4745__A _4855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3960_ _5725_/Q _3983_/B vssd1 vssd1 vccd1 vccd1 _3960_/Y sky130_fd_sc_hd__nand2_1
XFILLER_35_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2911_ _3844_/C vssd1 vssd1 vccd1 vccd1 _3288_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_50_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3891_ _3891_/A _3891_/B vssd1 vssd1 vccd1 vccd1 _3891_/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2842_ _5327_/A _5309_/A _5297_/A vssd1 vssd1 vccd1 vccd1 _3063_/C sky130_fd_sc_hd__nor3_1
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5630_ _5353_/X _5623_/X _5629_/X _5627_/X vssd1 vssd1 vccd1 vccd1 _6114_/D sky130_fd_sc_hd__o211a_1
X_5561_ _5577_/B vssd1 vssd1 vccd1 vccd1 _5570_/B sky130_fd_sc_hd__clkbuf_1
X_4512_ _5284_/A _4512_/B _4514_/B vssd1 vssd1 vccd1 vccd1 _5861_/D sky130_fd_sc_hd__nor3_1
XANTENNA__3096__A _3928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5492_ _5535_/B _5622_/B vssd1 vssd1 vccd1 vccd1 _5493_/A sky130_fd_sc_hd__or2_1
X_4443_ _3111_/X _4442_/X _3886_/A vssd1 vssd1 vccd1 vccd1 _4443_/X sky130_fd_sc_hd__o21a_1
XANTENNA__3824__A _3824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4374_ _5828_/Q _4373_/X _4374_/S vssd1 vssd1 vccd1 vccd1 _4375_/A sky130_fd_sc_hd__mux2_1
X_3325_ _3906_/B _3484_/A vssd1 vssd1 vccd1 vccd1 _3483_/A sky130_fd_sc_hd__or2_1
XFILLER_58_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6113_ _6115_/CLK _6113_/D vssd1 vssd1 vccd1 vccd1 _6113_/Q sky130_fd_sc_hd__dfxtp_1
X_3256_ _3256_/A vssd1 vssd1 vccd1 vccd1 _3522_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6044_ _6117_/CLK _6044_/D vssd1 vssd1 vccd1 vccd1 _6044_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3112__A1 _3820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3187_ _5910_/Q vssd1 vssd1 vccd1 vccd1 _4928_/A sky130_fd_sc_hd__inv_2
XANTENNA__4655__A _4914_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_383 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4612__A1 _5667_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5828_ _6101_/CLK _5828_/D vssd1 vssd1 vccd1 vccd1 _5828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5759_ _5777_/CLK _5759_/D vssd1 vssd1 vccd1 vccd1 _5759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4128__A0 _6118_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5325__C1 _3867_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_139 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3406__A2 _3484_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4603__A1 _6041_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3878__C1 _4210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3110_ _3282_/B vssd1 vssd1 vccd1 vccd1 _3821_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4090_ _5770_/Q _4089_/X _4097_/S vssd1 vssd1 vccd1 vccd1 _4091_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3041_ _3874_/A _3045_/B vssd1 vssd1 vccd1 vccd1 _3042_/A sky130_fd_sc_hd__nor2_1
XFILLER_48_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_512 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4992_ _5929_/Q _4993_/C _4991_/Y vssd1 vssd1 vccd1 vccd1 _5929_/D sky130_fd_sc_hd__a21oi_1
XFILLER_90_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3943_ _3979_/A _3943_/B vssd1 vssd1 vccd1 vccd1 _5722_/D sky130_fd_sc_hd__nor2_1
X_3874_ _3874_/A _3874_/B _5229_/B vssd1 vssd1 vccd1 vccd1 _3874_/X sky130_fd_sc_hd__and3_1
XFILLER_31_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5613_ _3604_/X _5602_/X _5611_/X _5612_/X vssd1 vssd1 vccd1 vccd1 _6108_/D sky130_fd_sc_hd__o211a_1
XFILLER_8_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5544_ _5544_/A vssd1 vssd1 vccd1 vccd1 _5597_/A sky130_fd_sc_hd__clkbuf_2
X_5475_ _6058_/Q _5483_/B vssd1 vssd1 vccd1 vccd1 _5475_/X sky130_fd_sc_hd__or2_1
XANTENNA__3581__A1 _3563_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4426_ _5973_/Q _5843_/Q _4426_/S vssd1 vssd1 vccd1 vccd1 _4426_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4357_ _5823_/Q _4356_/X _4357_/S vssd1 vssd1 vccd1 vccd1 _4358_/A sky130_fd_sc_hd__mux2_1
Xuser_proj_example_94 vssd1 vssd1 vccd1 vccd1 user_proj_example_94/HI io_oeb[12] sky130_fd_sc_hd__conb_1
Xuser_proj_example_83 vssd1 vssd1 vccd1 vccd1 user_proj_example_83/HI io_oeb[0] sky130_fd_sc_hd__conb_1
X_3308_ _3841_/B vssd1 vssd1 vccd1 vccd1 _3466_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4288_ _4288_/A _4329_/B vssd1 vssd1 vccd1 vccd1 _4288_/Y sky130_fd_sc_hd__nor2_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6027_ _6027_/CLK _6027_/D vssd1 vssd1 vccd1 vccd1 _6027_/Q sky130_fd_sc_hd__dfxtp_1
X_3239_ _5401_/A _5933_/Q _5927_/Q _5384_/A _3238_/Y vssd1 vssd1 vccd1 vccd1 _3243_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_39_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3729__A _3732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_478 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4588__A0 _5713_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3590_ _3593_/A vssd1 vssd1 vccd1 vccd1 _5601_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__4760__A0 _5657_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5260_ _5260_/A _5260_/B _5259_/X _3929_/C vssd1 vssd1 vccd1 vccd1 _5261_/C sky130_fd_sc_hd__or4bb_1
X_4211_ _5241_/A _6123_/Q _3814_/B vssd1 vssd1 vccd1 vccd1 _4211_/X sky130_fd_sc_hd__a21o_1
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5191_ _5191_/A vssd1 vssd1 vccd1 vccd1 _5993_/D sky130_fd_sc_hd__clkbuf_1
X_4142_ _6135_/Q _5784_/Q _4145_/S vssd1 vssd1 vccd1 vccd1 _4142_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4917__B _4917_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3821__B _3891_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4073_ _5765_/Q _4072_/X _4080_/S vssd1 vssd1 vccd1 vccd1 _4074_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4409__S _4409_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3024_ _3839_/A vssd1 vssd1 vccd1 vccd1 _3853_/A sky130_fd_sc_hd__buf_2
XFILLER_55_139 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_13_wb_clk_i clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6012_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_36_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4975_ _5924_/Q _4975_/B vssd1 vssd1 vccd1 vccd1 _4975_/X sky130_fd_sc_hd__and2_1
XFILLER_51_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3926_ _4210_/A _3925_/Y _5745_/Q _5746_/Q vssd1 vssd1 vccd1 vccd1 _3930_/A sky130_fd_sc_hd__o211a_1
XFILLER_51_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3857_ _5721_/Q _3857_/B vssd1 vssd1 vccd1 vccd1 _5234_/B sky130_fd_sc_hd__nand2_2
X_3788_ _3614_/A _5711_/Q _3791_/S vssd1 vssd1 vccd1 vccd1 _3789_/B sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_25_wb_clk_i_A clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_3_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5527_ _5393_/X _5514_/X _5526_/X _5518_/X vssd1 vssd1 vccd1 vccd1 _6077_/D sky130_fd_sc_hd__o211a_1
XFILLER_3_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5458_ _6052_/Q _5460_/B vssd1 vssd1 vccd1 vccd1 _5458_/X sky130_fd_sc_hd__or2_1
XFILLER_59_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4409_ _6062_/Q _5838_/Q _4409_/S vssd1 vssd1 vccd1 vccd1 _4409_/X sky130_fd_sc_hd__mux2_1
X_5389_ _5389_/A vssd1 vssd1 vccd1 vccd1 _5389_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_86_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3459__A _5279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3545__A1 _3221_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3360__C _3821_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4760_ _5657_/Q _4759_/X _4770_/S vssd1 vssd1 vccd1 vccd1 _4760_/X sky130_fd_sc_hd__mux2_1
X_3711_ _3711_/A vssd1 vssd1 vccd1 vccd1 _4594_/A sky130_fd_sc_hd__inv_2
X_4691_ _5102_/A vssd1 vssd1 vccd1 vccd1 _4732_/B sky130_fd_sc_hd__clkbuf_1
X_3642_ _3648_/A _3642_/B vssd1 vssd1 vccd1 vccd1 _3643_/A sky130_fd_sc_hd__and2_1
X_5312_ _5315_/A _5315_/B _5281_/B _5244_/B vssd1 vssd1 vccd1 vccd1 _5312_/X sky130_fd_sc_hd__a31o_1
X_3573_ _5343_/A _3738_/A vssd1 vssd1 vccd1 vccd1 _3577_/A sky130_fd_sc_hd__nand2_1
XFILLER_5_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5243_ _5243_/A _5243_/B vssd1 vssd1 vccd1 vccd1 _5271_/B sky130_fd_sc_hd__nand2_1
X_5174_ _5174_/A _5201_/B vssd1 vssd1 vccd1 vccd1 _5198_/S sky130_fd_sc_hd__nand2_2
XANTENNA__3551__B _5713_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4125_ _6117_/Q _5779_/Q _4128_/S vssd1 vssd1 vccd1 vccd1 _4125_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4056_ _5760_/Q _4055_/X _4063_/S vssd1 vssd1 vccd1 vccd1 _4057_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3007_ _3824_/D _3484_/A _3007_/C vssd1 vssd1 vccd1 vccd1 _3007_/X sky130_fd_sc_hd__or3_1
XFILLER_64_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4958_ _5920_/Q _4958_/B vssd1 vssd1 vccd1 vccd1 _4959_/B sky130_fd_sc_hd__xnor2_1
XFILLER_51_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3909_ _3917_/A _3875_/X _3908_/X _4554_/S vssd1 vssd1 vccd1 vccd1 _3909_/X sky130_fd_sc_hd__o211a_1
X_4889_ _5904_/Q _4858_/X _4887_/X _4888_/X vssd1 vssd1 vccd1 vccd1 _5904_/D sky130_fd_sc_hd__a22o_1
XANTENNA__5494__A _5537_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_286 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_426 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4246__A2 _4228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5579__A _5579_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5930_ _5959_/CLK _5930_/D vssd1 vssd1 vccd1 vccd1 _5930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5861_ _5926_/CLK _5861_/D vssd1 vssd1 vccd1 vccd1 _5861_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3099__A _4210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4812_ _6109_/Q _4811_/X _4822_/S vssd1 vssd1 vccd1 vccd1 _4812_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5792_ _6109_/CLK _5792_/D vssd1 vssd1 vccd1 vccd1 _5792_/Q sky130_fd_sc_hd__dfxtp_1
X_4743_ _6054_/Q _4706_/X _4716_/X _4742_/X vssd1 vssd1 vccd1 vccd1 _4743_/X sky130_fd_sc_hd__a211o_1
X_4674_ _5403_/B vssd1 vssd1 vccd1 vccd1 _4674_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3625_ _3794_/A _4645_/S vssd1 vssd1 vccd1 vccd1 _5174_/A sky130_fd_sc_hd__and2_2
X_3556_ _3556_/A _3556_/B vssd1 vssd1 vccd1 vccd1 _3556_/Y sky130_fd_sc_hd__nor2_1
XFILLER_88_326 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3487_ _3483_/A _3480_/X _3483_/X _3484_/X _3486_/X vssd1 vssd1 vccd1 vccd1 _3487_/X
+ sky130_fd_sc_hd__o2111a_1
X_5226_ _5295_/A _5226_/B vssd1 vssd1 vccd1 vccd1 _5227_/A sky130_fd_sc_hd__and2_1
X_5157_ _5408_/A vssd1 vssd1 vccd1 vccd1 _5391_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_29_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4108_ _5775_/Q _4107_/X _4116_/S vssd1 vssd1 vccd1 vccd1 _4109_/A sky130_fd_sc_hd__mux2_1
X_5088_ _5056_/X _5080_/X _5085_/X _5087_/X vssd1 vssd1 vccd1 vccd1 _5956_/D sky130_fd_sc_hd__o211a_1
XANTENNA__2906__A _3824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4039_ _5755_/Q _4038_/X _4046_/S vssd1 vssd1 vccd1 vccd1 _4040_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_462 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3920__A1 _6120_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input35_A la_data_in[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5399__A _6031_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_proj_example_120 vssd1 vssd1 vccd1 vccd1 user_proj_example_120/HI io_out[1]
+ sky130_fd_sc_hd__conb_1
XFILLER_11_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_proj_example_153 vssd1 vssd1 vccd1 vccd1 user_proj_example_153/HI la_data_out[28]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_131 vssd1 vssd1 vccd1 vccd1 user_proj_example_131/HI la_data_out[6]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_142 vssd1 vssd1 vccd1 vccd1 user_proj_example_142/HI la_data_out[17]
+ sky130_fd_sc_hd__conb_1
X_3410_ _3410_/A _3466_/D _3410_/C vssd1 vssd1 vccd1 vccd1 _3410_/X sky130_fd_sc_hd__and3_1
XFILLER_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_proj_example_186 vssd1 vssd1 vccd1 vccd1 user_proj_example_186/HI la_data_out[61]
+ sky130_fd_sc_hd__conb_1
X_4390_ _6055_/Q _5832_/Q _4396_/S vssd1 vssd1 vccd1 vccd1 _4390_/X sky130_fd_sc_hd__mux2_1
Xuser_proj_example_164 vssd1 vssd1 vccd1 vccd1 user_proj_example_164/HI la_data_out[39]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_175 vssd1 vssd1 vccd1 vccd1 user_proj_example_175/HI la_data_out[50]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_197 vssd1 vssd1 vccd1 vccd1 user_proj_example_197/HI la_data_out[104]
+ sky130_fd_sc_hd__conb_1
X_3341_ _3350_/C _3341_/B vssd1 vssd1 vccd1 vccd1 _4239_/B sky130_fd_sc_hd__nor2_1
XANTENNA__5581__B _5601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3272_ _4436_/A _3272_/B vssd1 vssd1 vccd1 vccd1 _3272_/Y sky130_fd_sc_hd__nor2_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6060_ _6108_/CLK _6060_/D vssd1 vssd1 vccd1 vccd1 _6060_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_510 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5011_ _5011_/A _5011_/B vssd1 vssd1 vccd1 vccd1 _5025_/B sky130_fd_sc_hd__nor2_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5416__A1 _3604_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5913_ _5920_/CLK _5913_/D vssd1 vssd1 vccd1 vccd1 _5913_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5844_ _5944_/CLK _5844_/D vssd1 vssd1 vccd1 vccd1 _5844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2987_ _3841_/A _3837_/A vssd1 vssd1 vccd1 vccd1 _3116_/A sky130_fd_sc_hd__nand2_1
X_5775_ _5941_/CLK _5775_/D vssd1 vssd1 vccd1 vccd1 _5775_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4152__S _4162_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4726_ _5888_/Q _4705_/X _4724_/X _4725_/X vssd1 vssd1 vccd1 vccd1 _5888_/D sky130_fd_sc_hd__a22o_1
X_4657_ _6118_/Q _4656_/X _4667_/S vssd1 vssd1 vccd1 vccd1 _4657_/X sky130_fd_sc_hd__mux2_1
X_3608_ _5662_/Q _3608_/B vssd1 vssd1 vccd1 vccd1 _3608_/X sky130_fd_sc_hd__or2_1
X_4588_ _5713_/Q _5666_/Q _4914_/S vssd1 vssd1 vccd1 vccd1 _4588_/X sky130_fd_sc_hd__mux2_1
X_3539_ _4548_/A _3537_/X _3538_/Y vssd1 vssd1 vccd1 vccd1 _3544_/C sky130_fd_sc_hd__o21a_1
XFILLER_88_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3723__C _3723_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5655__A1 _5396_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5209_ _5209_/A vssd1 vssd1 vccd1 vccd1 _5998_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4449__A2 _3331_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3930__A _3930_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3121__A2 _3938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2910_ _2949_/C _2949_/D vssd1 vssd1 vccd1 vccd1 _3844_/C sky130_fd_sc_hd__nor2_1
XFILLER_50_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3890_ _3890_/A vssd1 vssd1 vccd1 vccd1 _5718_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2841_ _6010_/Q vssd1 vssd1 vccd1 vccd1 _5297_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5560_ _5603_/B _5624_/B vssd1 vssd1 vccd1 vccd1 _5577_/B sky130_fd_sc_hd__nor2_1
X_4511_ _4511_/A _4511_/B vssd1 vssd1 vccd1 vccd1 _4514_/B sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_38_wb_clk_i clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5974_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_5491_ _3617_/X _5470_/A _5490_/X _5488_/X vssd1 vssd1 vccd1 vccd1 _6064_/D sky130_fd_sc_hd__o211a_1
X_4442_ _3867_/A _4437_/Y _4441_/X _3435_/A vssd1 vssd1 vccd1 vccd1 _4442_/X sky130_fd_sc_hd__o31a_1
XANTENNA__5592__A _6101_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3824__B _4002_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4373_ _6050_/Q _5827_/Q _4380_/S vssd1 vssd1 vccd1 vccd1 _4373_/X sky130_fd_sc_hd__mux2_1
X_3324_ _3896_/A _4466_/B vssd1 vssd1 vccd1 vccd1 _3906_/B sky130_fd_sc_hd__nand2_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6112_ _6112_/CLK _6112_/D vssd1 vssd1 vccd1 vccd1 _6112_/Q sky130_fd_sc_hd__dfxtp_1
X_3255_ _3668_/A vssd1 vssd1 vccd1 vccd1 _3255_/X sky130_fd_sc_hd__clkbuf_2
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6043_ _6117_/CLK _6043_/D vssd1 vssd1 vccd1 vccd1 _6043_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3840__A _4002_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3186_ _3186_/A _5916_/Q vssd1 vssd1 vccd1 vccd1 _3186_/Y sky130_fd_sc_hd__nor2_1
XFILLER_54_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5827_ _6101_/CLK _5827_/D vssd1 vssd1 vccd1 vccd1 _5827_/Q sky130_fd_sc_hd__dfxtp_1
X_5758_ _6005_/CLK _5758_/D vssd1 vssd1 vccd1 vccd1 _5758_/Q sky130_fd_sc_hd__dfxtp_1
X_4709_ _6135_/Q _4708_/X _4719_/S vssd1 vssd1 vccd1 vccd1 _4709_/X sky130_fd_sc_hd__mux2_1
X_5689_ _5996_/CLK _5689_/D vssd1 vssd1 vccd1 vccd1 _5689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5628__A1 _5342_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3750__A _3750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3811__B1 _3525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5619__A1 _3614_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3040_ _3463_/B _3040_/B vssd1 vssd1 vccd1 vccd1 _3045_/B sky130_fd_sc_hd__and2_1
XFILLER_36_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4055__A0 _6102_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4991_ _5929_/Q _4993_/C _4990_/X vssd1 vssd1 vccd1 vccd1 _4991_/Y sky130_fd_sc_hd__o21ai_1
X_3942_ _5722_/Q _3932_/X _3941_/X vssd1 vssd1 vccd1 vccd1 _3943_/B sky130_fd_sc_hd__a21oi_1
XFILLER_16_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3873_ _3873_/A _3873_/B _3873_/C _3873_/D vssd1 vssd1 vccd1 vccd1 _5229_/B sky130_fd_sc_hd__or4_1
X_5612_ _5638_/A vssd1 vssd1 vccd1 vccd1 _5612_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5543_ _6083_/Q _5549_/B vssd1 vssd1 vccd1 vccd1 _5543_/X sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_15_wb_clk_i_A clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_5474_ _3587_/X _5470_/X _5473_/X _5461_/X vssd1 vssd1 vccd1 vccd1 _6057_/D sky130_fd_sc_hd__o211a_1
X_4425_ _4425_/A vssd1 vssd1 vccd1 vccd1 _5843_/D sky130_fd_sc_hd__clkbuf_1
X_4356_ _6045_/Q _5822_/Q _4363_/S vssd1 vssd1 vccd1 vccd1 _4356_/X sky130_fd_sc_hd__mux2_1
X_3307_ _3460_/A _3857_/B _4550_/A vssd1 vssd1 vccd1 vccd1 _3462_/C sky130_fd_sc_hd__or3_1
XFILLER_58_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_proj_example_95 vssd1 vssd1 vccd1 vccd1 user_proj_example_95/HI io_oeb[13] sky130_fd_sc_hd__conb_1
Xuser_proj_example_84 vssd1 vssd1 vccd1 vccd1 user_proj_example_84/HI io_oeb[2] sky130_fd_sc_hd__conb_1
XFILLER_86_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4287_ _4287_/A _4287_/B vssd1 vssd1 vccd1 vccd1 _4291_/C sky130_fd_sc_hd__nand2_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6026_ _6027_/CLK _6026_/D vssd1 vssd1 vccd1 vccd1 _6026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3238_ _6030_/Q _5931_/Q vssd1 vssd1 vccd1 vccd1 _3238_/Y sky130_fd_sc_hd__xnor2_1
X_3169_ _4322_/A _3522_/A _3484_/B _3167_/X _3350_/A vssd1 vssd1 vccd1 vccd1 _3170_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_66_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5491__C1 _5488_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_54_wb_clk_i_A clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_10_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3021__A1 _3375_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_479 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3480__A _3480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4588__A1 _5666_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4210_ _4210_/A _4210_/B vssd1 vssd1 vccd1 vccd1 _4210_/Y sky130_fd_sc_hd__nor2_1
XFILLER_5_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5190_ _5204_/A _5190_/B vssd1 vssd1 vccd1 vccd1 _5191_/A sky130_fd_sc_hd__and2_1
X_4141_ _4141_/A vssd1 vssd1 vccd1 vccd1 _5784_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3821__C _3821_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4072_ _6108_/Q _5764_/Q _4075_/S vssd1 vssd1 vccd1 vccd1 _4072_/X sky130_fd_sc_hd__mux2_1
X_3023_ _4280_/A vssd1 vssd1 vccd1 vccd1 _3839_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4974_ _5924_/Q _4955_/X _4972_/X _4973_/Y _5284_/A vssd1 vssd1 vccd1 vccd1 _5924_/D
+ sky130_fd_sc_hd__a311oi_1
XFILLER_63_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3925_ _5747_/Q vssd1 vssd1 vccd1 vccd1 _3925_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_53_wb_clk_i clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6031_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3856_ _3913_/A _5233_/C vssd1 vssd1 vccd1 vccd1 _4010_/A sky130_fd_sc_hd__or2_1
XANTENNA__3408__C_N _4366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3787_ _5188_/A vssd1 vssd1 vccd1 vccd1 _3966_/A sky130_fd_sc_hd__clkbuf_4
X_5526_ _6077_/Q _5526_/B vssd1 vssd1 vccd1 vccd1 _5526_/X sky130_fd_sc_hd__or2_1
XANTENNA__4160__S _4167_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5457_ _5386_/X _5449_/X _5456_/X _5446_/X vssd1 vssd1 vccd1 vccd1 _6051_/D sky130_fd_sc_hd__o211a_1
X_4408_ _4408_/A vssd1 vssd1 vccd1 vccd1 _5838_/D sky130_fd_sc_hd__clkbuf_1
X_5388_ _5386_/X _5378_/X _5387_/Y _5371_/X vssd1 vssd1 vccd1 vccd1 _6027_/D sky130_fd_sc_hd__o211a_1
XFILLER_59_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4339_ _6069_/Q _3275_/X _4399_/S vssd1 vssd1 vccd1 vccd1 _4340_/A sky130_fd_sc_hd__mux2_1
X_6009_ _6132_/CLK _6009_/D vssd1 vssd1 vccd1 vccd1 _6009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5464__C1 _5461_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4843__B _4885_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3242__A1 _5387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3242__B2 _5384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4258__B1 _4259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_376 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3710_ _5876_/Q vssd1 vssd1 vccd1 vccd1 _4575_/A sky130_fd_sc_hd__inv_2
XFILLER_60_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4690_ _6097_/Q _4689_/X _4720_/S vssd1 vssd1 vccd1 vccd1 _4690_/X sky130_fd_sc_hd__mux2_1
X_3641_ input9/X _5670_/Q _3641_/S vssd1 vssd1 vccd1 vccd1 _3642_/B sky130_fd_sc_hd__mux2_1
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3572_ _5046_/A _5046_/B _3572_/C vssd1 vssd1 vccd1 vccd1 _3738_/A sky130_fd_sc_hd__and3_1
X_5311_ _5315_/B _5281_/B _5315_/A vssd1 vssd1 vccd1 vccd1 _5311_/Y sky130_fd_sc_hd__a21oi_1
X_5242_ _5243_/A _5304_/A _5245_/B vssd1 vssd1 vccd1 vccd1 _5244_/A sky130_fd_sc_hd__o21a_1
X_5173_ _4480_/A _4981_/B _3418_/Y _5012_/B _5172_/X vssd1 vssd1 vccd1 vccd1 _5988_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_68_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4124_ _4124_/A vssd1 vssd1 vccd1 vccd1 _5779_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5105__A _5537_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput1 io_in[1] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4206__C_N _3379_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4055_ _6102_/Q _5759_/Q _4058_/S vssd1 vssd1 vccd1 vccd1 _4055_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3006_ _5720_/Q _3849_/B vssd1 vssd1 vccd1 vccd1 _3007_/C sky130_fd_sc_hd__nand2_1
XFILLER_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4957_ _4957_/A _4958_/B _4966_/A vssd1 vssd1 vccd1 vccd1 _5919_/D sky130_fd_sc_hd__nor3_1
X_3908_ _3897_/B _4259_/A _3899_/A _3907_/X vssd1 vssd1 vccd1 vccd1 _3908_/X sky130_fd_sc_hd__o31a_1
X_4888_ _5982_/Q _4854_/X _4855_/X vssd1 vssd1 vccd1 vccd1 _4888_/X sky130_fd_sc_hd__o21a_1
X_3839_ _3839_/A _3839_/B _3839_/C _3839_/D vssd1 vssd1 vccd1 vccd1 _4555_/C sky130_fd_sc_hd__and4_1
X_5509_ _6071_/Q _5511_/B vssd1 vssd1 vccd1 vccd1 _5509_/X sky130_fd_sc_hd__or2_1
XFILLER_86_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4854__A _5403_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4715__A1 _5887_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5579__B _5601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5860_ _5926_/CLK _5860_/D vssd1 vssd1 vccd1 vccd1 _5860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4811_ _5662_/Q _4810_/X _4821_/S vssd1 vssd1 vccd1 vccd1 _4811_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5600__C1 _5597_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5791_ _6109_/CLK _5791_/D vssd1 vssd1 vccd1 vccd1 _5791_/Q sky130_fd_sc_hd__dfxtp_1
X_4742_ _4717_/X _4739_/X _4741_/X _4722_/X vssd1 vssd1 vccd1 vccd1 _4742_/X sky130_fd_sc_hd__o211a_1
X_4673_ _5345_/A vssd1 vssd1 vccd1 vccd1 _5403_/B sky130_fd_sc_hd__buf_2
X_3624_ _4860_/A vssd1 vssd1 vccd1 vccd1 _4645_/S sky130_fd_sc_hd__clkbuf_2
X_3555_ _5849_/Q _5804_/Q _3147_/B vssd1 vssd1 vccd1 vccd1 _3556_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__3843__A _4002_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3486_ _3486_/A _3486_/B _3485_/X vssd1 vssd1 vccd1 vccd1 _3486_/X sky130_fd_sc_hd__or3b_1
XFILLER_88_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5225_ _5075_/A _6004_/Q _5225_/S vssd1 vssd1 vccd1 vccd1 _5226_/B sky130_fd_sc_hd__mux2_1
XANTENNA__5131__A1 _5045_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5156_ _5981_/Q _5162_/B vssd1 vssd1 vccd1 vccd1 _5156_/X sky130_fd_sc_hd__or2_1
X_4107_ _5961_/Q _5774_/Q _4110_/S vssd1 vssd1 vccd1 vccd1 _4107_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4674__A _5403_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5087_ _5141_/A vssd1 vssd1 vccd1 vccd1 _5087_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3445__A1 _2955_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4038_ _6097_/Q _3491_/X _3821_/C vssd1 vssd1 vccd1 vccd1 _4038_/X sky130_fd_sc_hd__o21ba_1
XFILLER_37_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5989_ _6002_/CLK _5989_/D vssd1 vssd1 vccd1 vccd1 _5989_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4945__A1 _5981_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4613__S _5624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3920__A2 _3491_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input28_A la_data_in[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4584__A _4706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3928__A _3928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4936__A1 _6039_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xuser_proj_example_110 vssd1 vssd1 vccd1 vccd1 user_proj_example_110/HI io_oeb[28]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_121 vssd1 vssd1 vccd1 vccd1 user_proj_example_121/HI io_out[37]
+ sky130_fd_sc_hd__conb_1
XFILLER_11_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xuser_proj_example_132 vssd1 vssd1 vccd1 vccd1 user_proj_example_132/HI la_data_out[7]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_143 vssd1 vssd1 vccd1 vccd1 user_proj_example_143/HI la_data_out[18]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_154 vssd1 vssd1 vccd1 vccd1 user_proj_example_154/HI la_data_out[29]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_187 vssd1 vssd1 vccd1 vccd1 user_proj_example_187/HI la_data_out[62]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_165 vssd1 vssd1 vccd1 vccd1 user_proj_example_165/HI la_data_out[40]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_176 vssd1 vssd1 vccd1 vccd1 user_proj_example_176/HI la_data_out[51]
+ sky130_fd_sc_hd__conb_1
XANTENNA__3372__B1 _3469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3340_ _4220_/A _6123_/Q _5258_/A _4293_/A _4447_/A vssd1 vssd1 vccd1 vccd1 _3340_/X
+ sky130_fd_sc_hd__a221o_1
Xuser_proj_example_198 vssd1 vssd1 vccd1 vccd1 user_proj_example_198/HI la_data_out[105]
+ sky130_fd_sc_hd__conb_1
XANTENNA__5649__C1 _5172_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ _3161_/X _3274_/B _3261_/X _3263_/X _3270_/X vssd1 vssd1 vccd1 vccd1 _3271_/X
+ sky130_fd_sc_hd__a311o_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _5935_/Q _5008_/A _5009_/Y vssd1 vssd1 vccd1 vccd1 _5935_/D sky130_fd_sc_hd__o21a_1
XFILLER_87_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4467__A3 _4322_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4624__B1 _4623_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5912_ _5914_/CLK _5912_/D vssd1 vssd1 vccd1 vccd1 _5912_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5843_ _5959_/CLK _5843_/D vssd1 vssd1 vccd1 vccd1 _5843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2986_ _3049_/A vssd1 vssd1 vccd1 vccd1 _3841_/A sky130_fd_sc_hd__buf_2
X_5774_ _5944_/CLK _5774_/D vssd1 vssd1 vccd1 vccd1 _5774_/Q sky130_fd_sc_hd__dfxtp_1
X_4725_ _6028_/Q _4674_/X _4675_/X vssd1 vssd1 vccd1 vccd1 _4725_/X sky130_fd_sc_hd__o21a_1
X_4656_ _5694_/Q _5671_/Q _4697_/S vssd1 vssd1 vccd1 vccd1 _4656_/X sky130_fd_sc_hd__mux2_1
X_3607_ _3607_/A vssd1 vssd1 vccd1 vccd1 _3607_/X sky130_fd_sc_hd__clkbuf_2
X_4587_ _4860_/A vssd1 vssd1 vccd1 vccd1 _4914_/S sky130_fd_sc_hd__buf_2
XANTENNA__5352__A1 _5342_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3538_ _5859_/Q vssd1 vssd1 vccd1 vccd1 _3538_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4560__C1 _4460_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3469_ _3469_/A _3469_/B _3469_/C vssd1 vssd1 vccd1 vccd1 _3469_/X sky130_fd_sc_hd__or3_1
X_5208_ _5220_/A _5208_/B vssd1 vssd1 vccd1 vccd1 _5209_/A sky130_fd_sc_hd__and2_1
X_5139_ _5065_/X _5125_/X _5138_/X _5130_/X vssd1 vssd1 vccd1 vccd1 _5975_/D sky130_fd_sc_hd__o211a_1
XFILLER_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_8_wb_clk_i _5813_/CLK vssd1 vssd1 vccd1 vccd1 _5777_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__4851__B _4885_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4918__A1 _4717_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5591__A1 _5389_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2840_ _6011_/Q vssd1 vssd1 vccd1 vccd1 _5309_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4510_ _4518_/C _5860_/Q _4504_/B vssd1 vssd1 vccd1 vccd1 _4511_/B sky130_fd_sc_hd__a21oi_1
X_5490_ _6064_/Q _5490_/B vssd1 vssd1 vccd1 vccd1 _5490_/X sky130_fd_sc_hd__or2_1
X_4441_ _3849_/B _4440_/Y _3007_/C _4437_/B vssd1 vssd1 vccd1 vccd1 _4441_/X sky130_fd_sc_hd__o211a_1
XANTENNA__3393__A _3632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4372_ _4372_/A vssd1 vssd1 vccd1 vccd1 _5827_/D sky130_fd_sc_hd__clkbuf_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6111_ _6112_/CLK _6111_/D vssd1 vssd1 vccd1 vccd1 _6111_/Q sky130_fd_sc_hd__dfxtp_1
X_3323_ _3438_/A _3322_/X _3439_/A vssd1 vssd1 vccd1 vccd1 _4466_/B sky130_fd_sc_hd__o21ai_2
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3254_ _4251_/A vssd1 vssd1 vccd1 vccd1 _3668_/A sky130_fd_sc_hd__buf_2
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6042_ _6115_/CLK _6042_/D vssd1 vssd1 vccd1 vccd1 _6042_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3185_ _5919_/Q vssd1 vssd1 vccd1 vccd1 _4953_/A sky130_fd_sc_hd__inv_2
XFILLER_81_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_44_wb_clk_i_A clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__4163__S _4167_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5826_ _6101_/CLK _5826_/D vssd1 vssd1 vccd1 vccd1 _5826_/Q sky130_fd_sc_hd__dfxtp_1
X_2969_ _4229_/A _2969_/B vssd1 vssd1 vccd1 vccd1 _3360_/B sky130_fd_sc_hd__and2b_1
X_5757_ _6005_/CLK _5757_/D vssd1 vssd1 vccd1 vccd1 _5757_/Q sky130_fd_sc_hd__dfxtp_1
X_4708_ _5699_/Q _5676_/Q _4748_/S vssd1 vssd1 vccd1 vccd1 _4708_/X sky130_fd_sc_hd__mux2_1
X_5688_ _6003_/CLK _5688_/D vssd1 vssd1 vccd1 vccd1 _5688_/Q sky130_fd_sc_hd__dfxtp_1
X_4639_ _5102_/A vssd1 vssd1 vccd1 vccd1 _4683_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_78_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3887__A1 _3459_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5316__A1 _3491_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3939__B_N _3930_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output59_A _5886_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4990_ _4995_/B vssd1 vssd1 vccd1 vccd1 _4990_/X sky130_fd_sc_hd__clkbuf_1
X_3941_ _3941_/A vssd1 vssd1 vccd1 vccd1 _3941_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3872_ _2917_/A _4550_/A _4550_/B _3327_/X _3328_/B vssd1 vssd1 vccd1 vccd1 _3872_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_31_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5611_ _6108_/Q _5614_/B vssd1 vssd1 vccd1 vccd1 _5611_/X sky130_fd_sc_hd__or2_1
X_5542_ _3598_/X _5536_/X _5541_/X _5529_/X vssd1 vssd1 vccd1 vccd1 _6082_/D sky130_fd_sc_hd__o211a_1
X_5473_ _6057_/Q _5483_/B vssd1 vssd1 vccd1 vccd1 _5473_/X sky130_fd_sc_hd__or2_1
X_4424_ _5843_/Q _4423_/X _4433_/S vssd1 vssd1 vccd1 vccd1 _4425_/A sky130_fd_sc_hd__mux2_1
X_4355_ _4355_/A vssd1 vssd1 vccd1 vccd1 _5822_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3851__A _5250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3306_ _4280_/A _5851_/Q vssd1 vssd1 vccd1 vccd1 _4550_/A sky130_fd_sc_hd__xor2_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_proj_example_96 vssd1 vssd1 vccd1 vccd1 user_proj_example_96/HI io_oeb[14] sky130_fd_sc_hd__conb_1
Xuser_proj_example_85 vssd1 vssd1 vccd1 vccd1 user_proj_example_85/HI io_oeb[3] sky130_fd_sc_hd__conb_1
XFILLER_86_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4286_ _3839_/B _4210_/B _4285_/X vssd1 vssd1 vccd1 vccd1 _4287_/B sky130_fd_sc_hd__o21ai_1
XFILLER_58_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6025_ _6027_/CLK _6025_/D vssd1 vssd1 vccd1 vccd1 _6025_/Q sky130_fd_sc_hd__dfxtp_1
X_3237_ _6026_/Q vssd1 vssd1 vccd1 vccd1 _5384_/A sky130_fd_sc_hd__clkinv_2
X_3168_ _6129_/Q vssd1 vssd1 vccd1 vccd1 _3350_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_clkbuf_leaf_0_wb_clk_i_A clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_39_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3099_ _4210_/A _3928_/B vssd1 vssd1 vccd1 vccd1 _3508_/C sky130_fd_sc_hd__or2_1
X_5809_ _5942_/CLK _5809_/D vssd1 vssd1 vccd1 vccd1 _5809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3557__B1 _3221_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3480__B _3480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input10_A la_data_in[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4592__A _4883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5170__C1 _5169_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4140_ _5784_/Q _4139_/X _4150_/S vssd1 vssd1 vccd1 vccd1 _4141_/A sky130_fd_sc_hd__mux2_1
X_4071_ _4071_/A vssd1 vssd1 vccd1 vccd1 _5764_/D sky130_fd_sc_hd__clkbuf_1
X_3022_ _3022_/A _3022_/B _3022_/C _3021_/X vssd1 vssd1 vccd1 vccd1 _3022_/X sky130_fd_sc_hd__or4b_1
XFILLER_55_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4973_ _4948_/X _4975_/B _5924_/Q vssd1 vssd1 vccd1 vccd1 _4973_/Y sky130_fd_sc_hd__a21oi_1
X_3924_ _4436_/A vssd1 vssd1 vccd1 vccd1 _3979_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3855_ _3901_/A _3901_/B _3913_/B _3854_/Y vssd1 vssd1 vccd1 vccd1 _5233_/C sky130_fd_sc_hd__a211o_1
X_3786_ _4251_/A vssd1 vssd1 vccd1 vccd1 _5188_/A sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_22_wb_clk_i clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5874_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_5525_ _5389_/X _5514_/X _5524_/X _5518_/X vssd1 vssd1 vccd1 vccd1 _6076_/D sky130_fd_sc_hd__o211a_1
X_5456_ _6051_/Q _5460_/B vssd1 vssd1 vccd1 vccd1 _5456_/X sky130_fd_sc_hd__or2_1
XFILLER_59_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4407_ _5838_/Q _4406_/X _4417_/S vssd1 vssd1 vccd1 vccd1 _4408_/A sky130_fd_sc_hd__mux2_1
X_5387_ _5387_/A _5387_/B vssd1 vssd1 vccd1 vccd1 _5387_/Y sky130_fd_sc_hd__nand2_1
XFILLER_86_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4338_ _4338_/A vssd1 vssd1 vccd1 vccd1 _5817_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_28 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4267__A1 _3938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4269_ _4329_/B _4269_/B _4269_/C _4269_/D vssd1 vssd1 vccd1 vccd1 _4270_/C sky130_fd_sc_hd__or4_1
XANTENNA_input2_A la_data_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6008_ _6132_/CLK _6008_/D vssd1 vssd1 vccd1 vccd1 _6008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5519__A1 _5376_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3491__A _4095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5207__A0 _5056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_130 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3640_ _3640_/A vssd1 vssd1 vccd1 vccd1 _5669_/D sky130_fd_sc_hd__clkbuf_1
X_3571_ _5667_/Q _3794_/A vssd1 vssd1 vccd1 vccd1 _5343_/A sky130_fd_sc_hd__and2_1
X_5310_ _5310_/A vssd1 vssd1 vccd1 vccd1 _5315_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5241_ _5241_/A _5241_/B _5241_/C vssd1 vssd1 vccd1 vccd1 _5245_/B sky130_fd_sc_hd__and3_1
X_5172_ _5638_/A vssd1 vssd1 vccd1 vccd1 _5172_/X sky130_fd_sc_hd__clkbuf_4
X_4123_ _5779_/Q _4122_/X _4133_/S vssd1 vssd1 vccd1 vccd1 _4124_/A sky130_fd_sc_hd__mux2_1
X_4054_ _4054_/A vssd1 vssd1 vccd1 vccd1 _5759_/D sky130_fd_sc_hd__clkbuf_1
Xinput2 la_data_in[0] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_2
XFILLER_28_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3005_ _3849_/A _3853_/C _3005_/C vssd1 vssd1 vccd1 vccd1 _3293_/A sky130_fd_sc_hd__or3_2
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4956_ _4982_/C _4955_/X _3723_/C vssd1 vssd1 vccd1 vccd1 _4966_/A sky130_fd_sc_hd__a21o_1
XFILLER_51_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3907_ _5255_/A _3901_/B _5775_/Q vssd1 vssd1 vccd1 vccd1 _3907_/X sky130_fd_sc_hd__a21o_1
X_4887_ _5974_/Q _4859_/X _4869_/X _4886_/X vssd1 vssd1 vccd1 vccd1 _4887_/X sky130_fd_sc_hd__a211o_1
XFILLER_20_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3838_ _3838_/A _4281_/A vssd1 vssd1 vccd1 vccd1 _3839_/D sky130_fd_sc_hd__nor2_1
XANTENNA__4171__S _4184_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3769_ _3769_/A vssd1 vssd1 vccd1 vccd1 _5705_/D sky130_fd_sc_hd__clkbuf_1
X_5508_ _5366_/X _5493_/A _5507_/X _5503_/X vssd1 vssd1 vccd1 vccd1 _6070_/D sky130_fd_sc_hd__o211a_1
XFILLER_10_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5439_ _6045_/Q _5439_/B vssd1 vssd1 vccd1 vccd1 _5439_/X sky130_fd_sc_hd__or2_1
XFILLER_86_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4346__S _5278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4870__A _4870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5206__A _5408_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4651__A1 _6021_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4810_ _5709_/Q _5686_/Q _4848_/S vssd1 vssd1 vccd1 vccd1 _4810_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5790_ _6024_/CLK _5790_/D vssd1 vssd1 vccd1 vccd1 _5790_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3396__A _5234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4741_ _6078_/Q _4783_/B vssd1 vssd1 vccd1 vccd1 _4741_/X sky130_fd_sc_hd__or2_1
XFILLER_14_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4672_ _6047_/Q _4654_/X _4664_/X _4671_/X vssd1 vssd1 vccd1 vccd1 _4672_/X sky130_fd_sc_hd__a211o_1
X_3623_ _3712_/B _4597_/A vssd1 vssd1 vccd1 vccd1 _4860_/A sky130_fd_sc_hd__nor2_2
X_3554_ _3135_/C _5742_/Q vssd1 vssd1 vccd1 vccd1 _4530_/A sky130_fd_sc_hd__and2b_1
XFILLER_88_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3485_ _5245_/A _2863_/X _3428_/B _3851_/C vssd1 vssd1 vccd1 vccd1 _3485_/X sky130_fd_sc_hd__a31o_1
XFILLER_69_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5224_ _5224_/A vssd1 vssd1 vccd1 vccd1 _6003_/D sky130_fd_sc_hd__clkbuf_1
X_5155_ _5056_/X _5149_/X _5154_/X _5141_/X vssd1 vssd1 vccd1 vccd1 _5980_/D sky130_fd_sc_hd__o211a_1
XFILLER_56_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4106_ _4106_/A vssd1 vssd1 vccd1 vccd1 _5774_/D sky130_fd_sc_hd__clkbuf_1
X_5086_ _5408_/A vssd1 vssd1 vccd1 vccd1 _5141_/A sky130_fd_sc_hd__clkbuf_1
X_4037_ _4037_/A vssd1 vssd1 vccd1 vccd1 _5754_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5988_ _5988_/CLK _5988_/D vssd1 vssd1 vccd1 vccd1 _5988_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4939_ _4939_/A _4944_/B vssd1 vssd1 vccd1 vccd1 _4939_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_203 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2832__B _2880_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xuser_proj_example_111 vssd1 vssd1 vccd1 vccd1 user_proj_example_111/HI io_oeb[29]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_100 vssd1 vssd1 vccd1 vccd1 user_proj_example_100/HI io_oeb[18]
+ sky130_fd_sc_hd__conb_1
XFILLER_7_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3944__A _3954_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_proj_example_122 vssd1 vssd1 vccd1 vccd1 user_proj_example_122/HI irq[0] sky130_fd_sc_hd__conb_1
Xuser_proj_example_133 vssd1 vssd1 vccd1 vccd1 user_proj_example_133/HI la_data_out[8]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_144 vssd1 vssd1 vccd1 vccd1 user_proj_example_144/HI la_data_out[19]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_188 vssd1 vssd1 vccd1 vccd1 user_proj_example_188/HI la_data_out[63]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_155 vssd1 vssd1 vccd1 vccd1 user_proj_example_155/HI la_data_out[30]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_166 vssd1 vssd1 vccd1 vccd1 user_proj_example_166/HI la_data_out[41]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_177 vssd1 vssd1 vccd1 vccd1 user_proj_example_177/HI la_data_out[52]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_199 vssd1 vssd1 vccd1 vccd1 user_proj_example_199/HI la_data_out[106]
+ sky130_fd_sc_hd__conb_1
X_3270_ _3266_/Y _3891_/B _3269_/X vssd1 vssd1 vccd1 vccd1 _3270_/X sky130_fd_sc_hd__a21o_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5911_ _5920_/CLK _5911_/D vssd1 vssd1 vccd1 vccd1 _5911_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4624__A1 _5354_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_34_wb_clk_i_A clkbuf_3_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_46_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5842_ _5929_/CLK _5842_/D vssd1 vssd1 vccd1 vccd1 _5842_/Q sky130_fd_sc_hd__dfxtp_1
X_5773_ _5944_/CLK _5773_/D vssd1 vssd1 vccd1 vccd1 _5773_/Q sky130_fd_sc_hd__dfxtp_1
X_2985_ _4217_/A _4218_/B vssd1 vssd1 vccd1 vccd1 _3435_/A sky130_fd_sc_hd__nand2_1
X_4724_ _6052_/Q _4706_/X _4716_/X _4723_/X vssd1 vssd1 vccd1 vccd1 _4724_/X sky130_fd_sc_hd__a211o_1
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3854__A _3854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4655_ _4914_/S vssd1 vssd1 vccd1 vccd1 _4697_/S sky130_fd_sc_hd__clkbuf_2
X_4586_ _4870_/A vssd1 vssd1 vccd1 vccd1 _4717_/A sky130_fd_sc_hd__clkbuf_2
X_3606_ _3604_/X _3592_/X _3605_/X _3585_/X vssd1 vssd1 vccd1 vccd1 _5661_/D sky130_fd_sc_hd__o211a_1
X_3537_ _4545_/B _4541_/A _4534_/A _4545_/A vssd1 vssd1 vccd1 vccd1 _3537_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3573__B _3738_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3468_ _3460_/X _3462_/X _3467_/Y _3483_/A vssd1 vssd1 vccd1 vccd1 _3468_/X sky130_fd_sc_hd__a31o_1
XFILLER_69_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3399_ _4241_/A vssd1 vssd1 vccd1 vccd1 _3802_/B sky130_fd_sc_hd__clkbuf_2
X_5207_ _5056_/A _5998_/Q _5216_/S vssd1 vssd1 vccd1 vccd1 _5208_/B sky130_fd_sc_hd__mux2_1
XFILLER_29_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5138_ _5975_/Q _5138_/B vssd1 vssd1 vccd1 vccd1 _5138_/X sky130_fd_sc_hd__or2_1
XFILLER_29_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5069_ _5069_/A vssd1 vssd1 vccd1 vccd1 _5069_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_44_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input40_A wb_rst_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4595__A _4842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5567__C1 _5556_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4440_ _4438_/X _4439_/X _5234_/B vssd1 vssd1 vccd1 vccd1 _4440_/Y sky130_fd_sc_hd__a21boi_1
X_4371_ _5827_/Q _4370_/X _4374_/S vssd1 vssd1 vccd1 vccd1 _4372_/A sky130_fd_sc_hd__mux2_1
X_6110_ _6112_/CLK _6110_/D vssd1 vssd1 vccd1 vccd1 _6110_/Q sky130_fd_sc_hd__dfxtp_1
X_3322_ _3322_/A vssd1 vssd1 vccd1 vccd1 _3322_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_3_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3253_ _5339_/S vssd1 vssd1 vccd1 vccd1 _5336_/S sky130_fd_sc_hd__clkbuf_2
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6041_ _6118_/CLK _6041_/D vssd1 vssd1 vccd1 vccd1 _6041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3184_ _3180_/Y _5917_/Q _5916_/Q _3186_/A _3183_/X vssd1 vssd1 vccd1 vccd1 _3196_/B
+ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_47_wb_clk_i clkbuf_3_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5996_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_534 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5825_ _6048_/CLK _5825_/D vssd1 vssd1 vccd1 vccd1 _5825_/Q sky130_fd_sc_hd__dfxtp_1
X_2968_ _5717_/Q _2997_/A vssd1 vssd1 vccd1 vccd1 _2969_/B sky130_fd_sc_hd__or2_1
X_5756_ _6005_/CLK _5756_/D vssd1 vssd1 vccd1 vccd1 _5756_/Q sky130_fd_sc_hd__dfxtp_1
X_4707_ _4914_/S vssd1 vssd1 vccd1 vccd1 _4748_/S sky130_fd_sc_hd__clkbuf_2
X_5687_ _5996_/CLK _5687_/D vssd1 vssd1 vccd1 vccd1 _5687_/Q sky130_fd_sc_hd__dfxtp_1
X_2899_ _2899_/A vssd1 vssd1 vccd1 vccd1 _3158_/A sky130_fd_sc_hd__clkbuf_2
X_4638_ _6092_/Q _4637_/X _4668_/S vssd1 vssd1 vccd1 vccd1 _4638_/X sky130_fd_sc_hd__mux2_1
X_4569_ _4567_/Y _3544_/B _3542_/A vssd1 vssd1 vccd1 vccd1 _4569_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_76_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_76 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3811__A2 _3379_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3327__A1 _3159_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4827__A1 _6038_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3940_ _3954_/B _3940_/B vssd1 vssd1 vccd1 vccd1 _3941_/A sky130_fd_sc_hd__nor2_1
XFILLER_63_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3871_ _3873_/A _3159_/B _2997_/A _3052_/A vssd1 vssd1 vccd1 vccd1 _4550_/B sky130_fd_sc_hd__o22a_1
XFILLER_83_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5610_ _3601_/X _5602_/X _5609_/X _5597_/X vssd1 vssd1 vccd1 vccd1 _6107_/D sky130_fd_sc_hd__o211a_1
X_5541_ _6082_/Q _5549_/B vssd1 vssd1 vccd1 vccd1 _5541_/X sky130_fd_sc_hd__or2_1
X_5472_ _5490_/B vssd1 vssd1 vccd1 vccd1 _5483_/B sky130_fd_sc_hd__clkbuf_1
X_4423_ _5972_/Q _5842_/Q _4426_/S vssd1 vssd1 vccd1 vccd1 _4423_/X sky130_fd_sc_hd__mux2_1
X_4354_ _5822_/Q _4353_/X _4357_/S vssd1 vssd1 vccd1 vccd1 _4355_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3305_ _3480_/A _3459_/D _2885_/B _3486_/B _3117_/B vssd1 vssd1 vccd1 vccd1 _3305_/X
+ sky130_fd_sc_hd__o32a_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_proj_example_86 vssd1 vssd1 vccd1 vccd1 user_proj_example_86/HI io_oeb[4] sky130_fd_sc_hd__conb_1
X_4285_ _5241_/A _5241_/C _3870_/A _3463_/B _3466_/C vssd1 vssd1 vccd1 vccd1 _4285_/X
+ sky130_fd_sc_hd__o32a_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5124__A _5469_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6024_ _6024_/CLK _6024_/D vssd1 vssd1 vccd1 vccd1 _6024_/Q sky130_fd_sc_hd__dfxtp_1
Xuser_proj_example_97 vssd1 vssd1 vccd1 vccd1 user_proj_example_97/HI io_oeb[15] sky130_fd_sc_hd__conb_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3236_ _6032_/Q vssd1 vssd1 vccd1 vccd1 _5401_/A sky130_fd_sc_hd__inv_2
XFILLER_39_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3167_ _3161_/X _3165_/X _4206_/A vssd1 vssd1 vccd1 vccd1 _3167_/X sky130_fd_sc_hd__a21o_1
X_3098_ _3481_/B _3118_/B _2852_/B _3159_/B vssd1 vssd1 vccd1 vccd1 _3928_/B sky130_fd_sc_hd__o22a_1
XANTENNA__4174__S _4184_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5808_ _5808_/CLK _5808_/D vssd1 vssd1 vccd1 vccd1 _5808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5739_ _6121_/CLK _5739_/D vssd1 vssd1 vccd1 vccd1 _5739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3309__A1 _5255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3480__C _3480_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_459 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5482__A1 _3604_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4113__A _4113_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4070_ _5764_/Q _4069_/X _4080_/S vssd1 vssd1 vccd1 vccd1 _4071_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3021_ _3375_/B _3841_/C _3016_/X _3019_/X _3046_/A vssd1 vssd1 vccd1 vccd1 _3021_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_36_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4972_ _4972_/A _4972_/B _4975_/B vssd1 vssd1 vccd1 vccd1 _4972_/X sky130_fd_sc_hd__or3_1
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3923_ _3923_/A vssd1 vssd1 vccd1 vccd1 _5721_/D sky130_fd_sc_hd__clkbuf_1
X_3854_ _3854_/A _3854_/B vssd1 vssd1 vccd1 vccd1 _3854_/Y sky130_fd_sc_hd__nor2_1
X_3785_ _3785_/A vssd1 vssd1 vccd1 vccd1 _5710_/D sky130_fd_sc_hd__clkbuf_1
X_5524_ _6076_/Q _5526_/B vssd1 vssd1 vccd1 vccd1 _5524_/X sky130_fd_sc_hd__or2_1
X_5455_ _5382_/X _5449_/X _5454_/X _5446_/X vssd1 vssd1 vccd1 vccd1 _6050_/D sky130_fd_sc_hd__o211a_1
X_4406_ _6061_/Q _5837_/Q _4409_/S vssd1 vssd1 vccd1 vccd1 _4406_/X sky130_fd_sc_hd__mux2_1
X_5386_ _5386_/A vssd1 vssd1 vccd1 vccd1 _5386_/X sky130_fd_sc_hd__buf_2
X_4337_ _6068_/Q _2944_/B _4337_/S vssd1 vssd1 vccd1 vccd1 _4338_/A sky130_fd_sc_hd__mux2_1
X_4268_ _3402_/Y _3459_/D _4233_/C vssd1 vssd1 vccd1 vccd1 _4269_/D sky130_fd_sc_hd__a21oi_1
X_6007_ _6012_/CLK _6007_/D vssd1 vssd1 vccd1 vccd1 _6007_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3219_ _3218_/X _5854_/Q vssd1 vssd1 vccd1 vccd1 _3219_/X sky130_fd_sc_hd__and2b_1
XANTENNA__4267__A2 _3480_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5464__A1 _5396_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4199_ _5952_/Q _5801_/Q _4554_/S vssd1 vssd1 vccd1 vccd1 _4199_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3102__A _4002_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3459__D _3459_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2941__A _2941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5455__A1 _5382_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_142 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3947__A _3966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2851__A _3049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3570_ _5987_/Q _3570_/B _3570_/C vssd1 vssd1 vccd1 vccd1 _3794_/A sky130_fd_sc_hd__and3b_2
X_5240_ _5240_/A _5257_/A vssd1 vssd1 vccd1 vccd1 _5287_/C sky130_fd_sc_hd__or2_1
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5171_ _5171_/A _5171_/B vssd1 vssd1 vccd1 vccd1 _5987_/D sky130_fd_sc_hd__nor2_1
XFILLER_68_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4122_ _6116_/Q _5778_/Q _4128_/S vssd1 vssd1 vccd1 vccd1 _4122_/X sky130_fd_sc_hd__mux2_1
X_4053_ _5759_/Q _4052_/X _4063_/S vssd1 vssd1 vccd1 vccd1 _4054_/A sky130_fd_sc_hd__mux2_1
X_3004_ _5720_/Q vssd1 vssd1 vccd1 vccd1 _3849_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput3 la_data_in[1] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_2
XFILLER_91_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_3_4__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4955_ _4964_/B vssd1 vssd1 vccd1 vccd1 _4955_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4452__S _4452_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3906_ _4210_/A _3906_/B vssd1 vssd1 vccd1 vccd1 _3917_/A sky130_fd_sc_hd__or2_1
X_4886_ _4870_/X _4884_/X _4885_/X _4875_/X vssd1 vssd1 vccd1 vccd1 _4886_/X sky130_fd_sc_hd__o211a_1
X_3837_ _3837_/A _3873_/D vssd1 vssd1 vccd1 vccd1 _3839_/C sky130_fd_sc_hd__nor2_1
X_3768_ _3768_/A _3768_/B vssd1 vssd1 vccd1 vccd1 _3769_/A sky130_fd_sc_hd__and2_1
X_5507_ _6070_/Q _5511_/B vssd1 vssd1 vccd1 vccd1 _5507_/X sky130_fd_sc_hd__or2_1
X_3699_ _3699_/A vssd1 vssd1 vccd1 vccd1 _5686_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5438_ _5360_/X _5427_/X _5437_/X _5435_/X vssd1 vssd1 vccd1 vccd1 _6044_/D sky130_fd_sc_hd__o211a_1
X_5369_ _5369_/A vssd1 vssd1 vccd1 vccd1 _5369_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_19_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4270__D_N _4228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_24_wb_clk_i_A clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_46_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5600__A1 _3582_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5061__C1 _5043_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4740_ _5102_/A vssd1 vssd1 vccd1 vccd1 _4783_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4671_ _4665_/X _4668_/X _4669_/X _4670_/X vssd1 vssd1 vccd1 vccd1 _4671_/X sky130_fd_sc_hd__o211a_1
X_3622_ _3711_/A _4591_/B vssd1 vssd1 vccd1 vccd1 _4597_/A sky130_fd_sc_hd__or2_1
X_3553_ _3553_/A _5742_/Q vssd1 vssd1 vccd1 vccd1 _3553_/X sky130_fd_sc_hd__and2_1
X_3484_ _3484_/A _3484_/B _3291_/C vssd1 vssd1 vccd1 vccd1 _3484_/X sky130_fd_sc_hd__or3b_1
X_5223_ _5295_/A _5223_/B vssd1 vssd1 vccd1 vccd1 _5224_/A sky130_fd_sc_hd__and2_1
X_5154_ _5980_/Q _5162_/B vssd1 vssd1 vccd1 vccd1 _5154_/X sky130_fd_sc_hd__or2_1
XFILLER_56_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4105_ _5774_/Q _4104_/X _4116_/S vssd1 vssd1 vccd1 vccd1 _4106_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5085_ _5956_/Q _5093_/B vssd1 vssd1 vccd1 vccd1 _5085_/X sky130_fd_sc_hd__or2_1
X_4036_ _5754_/Q _4035_/X _4046_/S vssd1 vssd1 vccd1 vccd1 _4037_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_443 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5987_ _6050_/CLK _5987_/D vssd1 vssd1 vccd1 vccd1 _5987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4938_ _6040_/Q _4928_/B _4937_/X _4929_/X vssd1 vssd1 vccd1 vccd1 _5914_/D sky130_fd_sc_hd__o211a_1
X_4869_ _4869_/A vssd1 vssd1 vccd1 vccd1 _4869_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4330__B2 _2955_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3497__A _5255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xuser_proj_example_112 vssd1 vssd1 vccd1 vccd1 user_proj_example_112/HI io_oeb[30]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_101 vssd1 vssd1 vccd1 vccd1 user_proj_example_101/HI io_oeb[19]
+ sky130_fd_sc_hd__conb_1
XFILLER_7_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_proj_example_123 vssd1 vssd1 vccd1 vccd1 user_proj_example_123/HI irq[1] sky130_fd_sc_hd__conb_1
Xuser_proj_example_134 vssd1 vssd1 vccd1 vccd1 user_proj_example_134/HI la_data_out[9]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_145 vssd1 vssd1 vccd1 vccd1 user_proj_example_145/HI la_data_out[20]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_178 vssd1 vssd1 vccd1 vccd1 user_proj_example_178/HI la_data_out[53]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_156 vssd1 vssd1 vccd1 vccd1 user_proj_example_156/HI la_data_out[31]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_167 vssd1 vssd1 vccd1 vccd1 user_proj_example_167/HI la_data_out[42]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_189 vssd1 vssd1 vccd1 vccd1 user_proj_example_189/HI la_data_out[96]
+ sky130_fd_sc_hd__conb_1
XANTENNA__5649__A1 _5386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4321__A1 _3494_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5910_ _5920_/CLK _5910_/D vssd1 vssd1 vccd1 vccd1 _5910_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4791__A _4842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5841_ _6040_/CLK _5841_/D vssd1 vssd1 vccd1 vccd1 _5841_/Q sky130_fd_sc_hd__dfxtp_1
X_2984_ _3300_/A _2983_/Y _3434_/A vssd1 vssd1 vccd1 vccd1 _2984_/X sky130_fd_sc_hd__o21a_1
X_5772_ _5914_/CLK _5772_/D vssd1 vssd1 vccd1 vccd1 _5772_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3200__A _6025_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4723_ _4717_/X _4720_/X _4721_/X _4722_/X vssd1 vssd1 vccd1 vccd1 _4723_/X sky130_fd_sc_hd__o211a_1
XANTENNA__3060__B2 _3272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4654_ _4706_/A vssd1 vssd1 vccd1 vccd1 _4654_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4585_ _4594_/A _4594_/B _4604_/B vssd1 vssd1 vccd1 vccd1 _4870_/A sky130_fd_sc_hd__nor3_2
X_3605_ _5661_/Q _3608_/B vssd1 vssd1 vccd1 vccd1 _3605_/X sky130_fd_sc_hd__or2_1
X_3536_ _5866_/Q vssd1 vssd1 vccd1 vccd1 _4534_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__5127__A _5471_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3467_ _3460_/C _3464_/Y _3466_/X vssd1 vssd1 vccd1 vccd1 _3467_/Y sky130_fd_sc_hd__a21oi_1
X_5206_ _5408_/A vssd1 vssd1 vccd1 vccd1 _5220_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_88_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3398_ _6124_/Q vssd1 vssd1 vccd1 vccd1 _4241_/A sky130_fd_sc_hd__inv_2
XFILLER_57_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4177__S _4184_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5137_ _5062_/X _5125_/X _5136_/X _5130_/X vssd1 vssd1 vccd1 vccd1 _5974_/D sky130_fd_sc_hd__o211a_1
XFILLER_72_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5068_ _5065_/X _5050_/X _5066_/X _5067_/X vssd1 vssd1 vccd1 vccd1 _5951_/D sky130_fd_sc_hd__o211a_1
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5273__C1 _4041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4019_ _5749_/Q _4018_/X _4028_/S vssd1 vssd1 vccd1 vccd1 _4020_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input33_A la_data_in[58] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5500__A _6067_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4370_ _6049_/Q _5826_/Q _4380_/S vssd1 vssd1 vccd1 vccd1 _4370_/X sky130_fd_sc_hd__mux2_1
X_3321_ _3321_/A vssd1 vssd1 vccd1 vccd1 _3438_/A sky130_fd_sc_hd__clkbuf_2
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3252_ _5240_/A vssd1 vssd1 vccd1 vccd1 _5339_/S sky130_fd_sc_hd__clkbuf_2
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6040_ _6040_/CLK _6040_/D vssd1 vssd1 vccd1 vccd1 _6040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3183_ _5920_/Q _4931_/A _4944_/A _5926_/Q vssd1 vssd1 vccd1 vccd1 _3183_/X sky130_fd_sc_hd__a2bb2o_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4058__A0 _6103_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_16_wb_clk_i _5836_/CLK vssd1 vssd1 vccd1 vccd1 _6018_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_34_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5824_ _6048_/CLK _5824_/D vssd1 vssd1 vccd1 vccd1 _5824_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_284 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2967_ _3859_/C vssd1 vssd1 vccd1 vccd1 _2997_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5755_ _6005_/CLK _5755_/D vssd1 vssd1 vccd1 vccd1 _5755_/Q sky130_fd_sc_hd__dfxtp_1
X_2898_ _3553_/A _3469_/A vssd1 vssd1 vccd1 vccd1 _2899_/A sky130_fd_sc_hd__nor2_1
X_5686_ _5996_/CLK _5686_/D vssd1 vssd1 vccd1 vccd1 _5686_/Q sky130_fd_sc_hd__dfxtp_1
X_4706_ _4706_/A vssd1 vssd1 vccd1 vccd1 _4706_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4637_ _6116_/Q _4636_/X _4667_/S vssd1 vssd1 vccd1 vccd1 _4637_/X sky130_fd_sc_hd__mux2_1
X_4568_ _5737_/Q _4568_/B vssd1 vssd1 vccd1 vccd1 _4568_/X sky130_fd_sc_hd__or2_1
XFILLER_1_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4499_ _5743_/Q _5740_/Q _5741_/Q vssd1 vssd1 vccd1 vccd1 _4501_/B sky130_fd_sc_hd__or3_1
X_3519_ _3405_/A _3516_/X _3517_/X _3518_/Y _3412_/A vssd1 vssd1 vccd1 vccd1 _3519_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_33 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3494__B _3494_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3870_ _3870_/A vssd1 vssd1 vccd1 vccd1 _5301_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_16_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5540_ _3587_/X _5536_/X _5539_/X _5529_/X vssd1 vssd1 vccd1 vccd1 _6081_/D sky130_fd_sc_hd__o211a_1
X_5471_ _5603_/A _5471_/B vssd1 vssd1 vccd1 vccd1 _5490_/B sky130_fd_sc_hd__nor2_1
XANTENNA__3318__A2 _3432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4422_ _4422_/A vssd1 vssd1 vccd1 vccd1 _5842_/D sky130_fd_sc_hd__clkbuf_1
X_4353_ _6044_/Q _5821_/Q _4363_/S vssd1 vssd1 vccd1 vccd1 _4353_/X sky130_fd_sc_hd__mux2_1
X_3304_ _3480_/B _3304_/B vssd1 vssd1 vccd1 vccd1 _3486_/B sky130_fd_sc_hd__nand2_1
X_4284_ _3480_/A _4279_/X _4282_/X _4283_/X vssd1 vssd1 vccd1 vccd1 _4291_/B sky130_fd_sc_hd__o211a_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_proj_example_87 vssd1 vssd1 vccd1 vccd1 user_proj_example_87/HI io_oeb[5] sky130_fd_sc_hd__conb_1
XFILLER_86_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6023_ _6024_/CLK _6023_/D vssd1 vssd1 vccd1 vccd1 _6023_/Q sky130_fd_sc_hd__dfxtp_2
X_3235_ _3230_/X _3231_/Y _3232_/Y _3233_/X _3234_/Y vssd1 vssd1 vccd1 vccd1 _3243_/B
+ sky130_fd_sc_hd__o221a_1
Xuser_proj_example_98 vssd1 vssd1 vccd1 vccd1 user_proj_example_98/HI io_oeb[16] sky130_fd_sc_hd__conb_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3166_ _3553_/A vssd1 vssd1 vccd1 vccd1 _4206_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_66_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3097_ _3814_/B vssd1 vssd1 vccd1 vccd1 _4210_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_54_335 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5140__A _5976_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_508 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4451__B1 _4449_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3298__C _3836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5807_ _6012_/CLK _5807_/D vssd1 vssd1 vccd1 vccd1 _5807_/Q sky130_fd_sc_hd__dfxtp_1
X_3999_ _3999_/A _3999_/B vssd1 vssd1 vccd1 vccd1 _5736_/D sky130_fd_sc_hd__nor2_1
XANTENNA__4203__A0 _5803_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5738_ _5874_/CLK _5738_/D vssd1 vssd1 vccd1 vccd1 _5738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4754__A1 _6031_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5669_ _6091_/CLK _5669_/D vssd1 vssd1 vccd1 vccd1 _5669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4690__A0 _6097_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2849__A _3038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output64_A _5891_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3020_ _3020_/A vssd1 vssd1 vccd1 vccd1 _3046_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_63_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4971_ _4971_/A vssd1 vssd1 vccd1 vccd1 _5923_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3922_ _3037_/A _3920_/X _3922_/S vssd1 vssd1 vccd1 vccd1 _3923_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3853_ _3853_/A _5720_/Q _3853_/C _3897_/D vssd1 vssd1 vccd1 vccd1 _3854_/B sky130_fd_sc_hd__or4_1
XANTENNA__4736__A1 _5889_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3784_ _3784_/A _3784_/B vssd1 vssd1 vccd1 vccd1 _3785_/A sky130_fd_sc_hd__and2_1
X_5523_ _5386_/X _5514_/X _5522_/X _5518_/X vssd1 vssd1 vccd1 vccd1 _6075_/D sky130_fd_sc_hd__o211a_1
X_5454_ _6050_/Q _5460_/B vssd1 vssd1 vccd1 vccd1 _5454_/X sky130_fd_sc_hd__or2_1
X_4405_ _6060_/Q _3802_/B _4417_/S _4404_/X vssd1 vssd1 vccd1 vccd1 _5837_/D sky130_fd_sc_hd__a31o_1
X_5385_ _5382_/X _5378_/X _5384_/Y _5371_/X vssd1 vssd1 vccd1 vccd1 _6026_/D sky130_fd_sc_hd__o211a_1
X_4336_ _4464_/B _4337_/S _4333_/Y _6067_/Q vssd1 vssd1 vccd1 vccd1 _5816_/D sky130_fd_sc_hd__a22o_1
XFILLER_59_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4267_ _3938_/A _3480_/C _4243_/A vssd1 vssd1 vccd1 vccd1 _4269_/C sky130_fd_sc_hd__o21a_1
XFILLER_59_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6006_ _6122_/CLK _6006_/D vssd1 vssd1 vccd1 vccd1 _6006_/Q sky130_fd_sc_hd__dfxtp_1
X_3218_ _4972_/A vssd1 vssd1 vccd1 vccd1 _3218_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_leaf_31_wb_clk_i _5836_/CLK vssd1 vssd1 vccd1 vccd1 _5941_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_39_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4198_ _4198_/A vssd1 vssd1 vccd1 vccd1 _5801_/D sky130_fd_sc_hd__clkbuf_1
X_3149_ _5859_/Q _5858_/Q _3546_/A _4480_/A vssd1 vssd1 vccd1 vccd1 _3149_/X sky130_fd_sc_hd__o31a_1
XANTENNA__3475__B2 _3480_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_18 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5301__C _5301_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5045__A _5045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_75 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_14_wb_clk_i_A clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_1_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_154 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2851__B _5736_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_53_wb_clk_i_A clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_5170_ _5075_/X _5149_/A _5168_/X _5169_/X vssd1 vssd1 vccd1 vccd1 _5986_/D sky130_fd_sc_hd__o211a_1
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4121_ _4121_/A vssd1 vssd1 vccd1 vccd1 _5778_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3457__A1 _3454_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4052_ _6101_/Q _5758_/Q _4058_/S vssd1 vssd1 vccd1 vccd1 _4052_/X sky130_fd_sc_hd__mux2_1
X_3003_ _3003_/A vssd1 vssd1 vccd1 vccd1 _3469_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_83_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput4 la_data_in[2] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3203__A _6024_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4954_ _4954_/A vssd1 vssd1 vccd1 vccd1 _4982_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3857__B _3857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3905_ _3905_/A vssd1 vssd1 vccd1 vccd1 _5719_/D sky130_fd_sc_hd__clkbuf_1
X_4885_ _5966_/Q _4885_/B vssd1 vssd1 vccd1 vccd1 _4885_/X sky130_fd_sc_hd__or2_1
X_3836_ _3836_/A _4288_/A vssd1 vssd1 vccd1 vccd1 _4555_/B sky130_fd_sc_hd__or2_1
X_3767_ _3587_/A _5705_/Q _3780_/S vssd1 vssd1 vccd1 vccd1 _3768_/B sky130_fd_sc_hd__mux2_1
XANTENNA__3873__A _3873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5506_ _5363_/X _5493_/X _5505_/X _5503_/X vssd1 vssd1 vccd1 vccd1 _6069_/D sky130_fd_sc_hd__o211a_1
X_3698_ _3701_/A _3698_/B vssd1 vssd1 vccd1 vccd1 _3699_/A sky130_fd_sc_hd__and2_1
XANTENNA__3145__A0 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5437_ _6044_/Q _5439_/B vssd1 vssd1 vccd1 vccd1 _5437_/X sky130_fd_sc_hd__or2_1
XFILLER_87_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5368_ _5366_/X _5354_/B _5367_/X _5355_/X vssd1 vssd1 vccd1 vccd1 _6022_/D sky130_fd_sc_hd__o211a_1
X_5299_ _5310_/A _5299_/B vssd1 vssd1 vccd1 vccd1 _5299_/Y sky130_fd_sc_hd__nor2_1
XFILLER_59_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4319_ _4016_/B _4318_/X _4014_/X vssd1 vssd1 vccd1 vccd1 _4319_/X sky130_fd_sc_hd__a21o_1
XANTENNA__2936__B _3317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3722__S _3722_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5503__A _5529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4636__A0 _5692_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4119__A _4170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2862__A _2941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4670_ _4824_/A vssd1 vssd1 vccd1 vccd1 _4670_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3621_ input3/X input2/X input4/X vssd1 vssd1 vccd1 vccd1 _4591_/B sky130_fd_sc_hd__or3b_1
X_3552_ _3550_/X _3551_/X _3245_/X vssd1 vssd1 vccd1 vccd1 _5741_/D sky130_fd_sc_hd__o21a_1
X_3483_ _3483_/A _3483_/B _3482_/Y vssd1 vssd1 vccd1 vccd1 _3483_/X sky130_fd_sc_hd__or3b_1
X_5222_ _5072_/A _6003_/Q _5225_/S vssd1 vssd1 vccd1 vccd1 _5223_/B sky130_fd_sc_hd__mux2_1
XFILLER_69_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5153_ _5045_/X _5149_/X _5152_/X _5141_/X vssd1 vssd1 vccd1 vccd1 _5979_/D sky130_fd_sc_hd__o211a_1
X_4104_ _5960_/Q _5773_/Q _4110_/S vssd1 vssd1 vccd1 vccd1 _4104_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5413__A _6035_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5084_ _5045_/X _5080_/X _5083_/X _5067_/X vssd1 vssd1 vccd1 vccd1 _5955_/D sky130_fd_sc_hd__o211a_1
XFILLER_56_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4035_ _6095_/Q _2858_/A _5753_/Q _4017_/A vssd1 vssd1 vccd1 vccd1 _4035_/X sky130_fd_sc_hd__a22o_1
XFILLER_2_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5986_ _5986_/CLK _5986_/D vssd1 vssd1 vccd1 vccd1 _5986_/Q sky130_fd_sc_hd__dfxtp_1
X_4937_ _5914_/Q _4942_/B vssd1 vssd1 vccd1 vccd1 _4937_/X sky130_fd_sc_hd__or2_1
X_4868_ _5902_/Q _4858_/X _4866_/X _4867_/X vssd1 vssd1 vccd1 vccd1 _5902_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3819_ _5336_/S _6016_/Q _4331_/B _3816_/B _3818_/X vssd1 vssd1 vccd1 vccd1 _5716_/D
+ sky130_fd_sc_hd__a41o_1
X_4799_ _6108_/Q _4798_/X _4822_/S vssd1 vssd1 vccd1 vccd1 _4799_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_proj_example_102 vssd1 vssd1 vccd1 vccd1 user_proj_example_102/HI io_oeb[20]
+ sky130_fd_sc_hd__conb_1
XFILLER_11_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_proj_example_113 vssd1 vssd1 vccd1 vccd1 user_proj_example_113/HI io_oeb[31]
+ sky130_fd_sc_hd__conb_1
XFILLER_7_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_proj_example_124 vssd1 vssd1 vccd1 vccd1 user_proj_example_124/HI irq[2] sky130_fd_sc_hd__conb_1
Xuser_proj_example_135 vssd1 vssd1 vccd1 vccd1 user_proj_example_135/HI la_data_out[10]
+ sky130_fd_sc_hd__conb_1
XFILLER_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_proj_example_168 vssd1 vssd1 vccd1 vccd1 user_proj_example_168/HI la_data_out[43]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_179 vssd1 vssd1 vccd1 vccd1 user_proj_example_179/HI la_data_out[54]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_146 vssd1 vssd1 vccd1 vccd1 user_proj_example_146/HI la_data_out[21]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_157 vssd1 vssd1 vccd1 vccd1 user_proj_example_157/HI la_data_out[32]
+ sky130_fd_sc_hd__conb_1
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5840_ _6112_/CLK _5840_/D vssd1 vssd1 vccd1 vccd1 _5840_/Q sky130_fd_sc_hd__dfxtp_1
X_2983_ _3020_/A _2983_/B vssd1 vssd1 vccd1 vccd1 _2983_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5771_ _5914_/CLK _5771_/D vssd1 vssd1 vccd1 vccd1 _5771_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4722_ _4824_/A vssd1 vssd1 vccd1 vccd1 _4722_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput40 wb_rst_i vssd1 vssd1 vccd1 vccd1 _2880_/A sky130_fd_sc_hd__clkbuf_2
X_4653_ _4756_/A vssd1 vssd1 vccd1 vccd1 _4653_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5408__A _5408_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3604_ _3604_/A vssd1 vssd1 vccd1 vccd1 _3604_/X sky130_fd_sc_hd__clkbuf_2
X_4584_ _4706_/A vssd1 vssd1 vccd1 vccd1 _4584_/X sky130_fd_sc_hd__clkbuf_2
X_3535_ _5867_/Q vssd1 vssd1 vccd1 vccd1 _4541_/A sky130_fd_sc_hd__clkbuf_1
X_3466_ _3466_/A _3840_/B _3466_/C _3466_/D vssd1 vssd1 vccd1 vccd1 _3466_/X sky130_fd_sc_hd__and4_1
X_5205_ _5205_/A vssd1 vssd1 vccd1 vccd1 _5997_/D sky130_fd_sc_hd__clkbuf_1
X_3397_ _4239_/B _3800_/B _3396_/Y _3117_/B vssd1 vssd1 vccd1 vccd1 _3397_/X sky130_fd_sc_hd__o211a_1
XFILLER_84_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5136_ _5974_/Q _5138_/B vssd1 vssd1 vccd1 vccd1 _5136_/X sky130_fd_sc_hd__or2_1
XFILLER_84_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5067_ _5067_/A vssd1 vssd1 vccd1 vccd1 _5067_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4018_ _6090_/Q _4014_/X _5748_/Q _4017_/X vssd1 vssd1 vccd1 vccd1 _4018_/X sky130_fd_sc_hd__a22o_1
XFILLER_25_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5969_ _5975_/CLK _5969_/D vssd1 vssd1 vccd1 vccd1 _5969_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5328__A1 _3491_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4303__A2 _3497_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input26_A la_data_in[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5264__B1 _3547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3290__A2 _3287_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5567__A1 _5357_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5228__A _5234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3320_ _3853_/C vssd1 vssd1 vccd1 vccd1 _3896_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3251_ _5256_/A vssd1 vssd1 vccd1 vccd1 _5240_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3182_ _5917_/Q vssd1 vssd1 vccd1 vccd1 _4944_/A sky130_fd_sc_hd__inv_2
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5823_ _6048_/CLK _5823_/D vssd1 vssd1 vccd1 vccd1 _5823_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2966_ _5808_/Q _5807_/Q _5806_/Q _5805_/Q vssd1 vssd1 vccd1 vccd1 _3859_/C sky130_fd_sc_hd__or4bb_1
XANTENNA__4230__A1 _5327_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5754_ _5796_/CLK _5754_/D vssd1 vssd1 vccd1 vccd1 _5754_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_56_wb_clk_i clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _5702_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2897_ _5279_/A vssd1 vssd1 vccd1 vccd1 _3469_/A sky130_fd_sc_hd__clkbuf_2
X_5685_ _6085_/CLK _5685_/D vssd1 vssd1 vccd1 vccd1 _5685_/Q sky130_fd_sc_hd__dfxtp_1
X_4705_ _4756_/A vssd1 vssd1 vccd1 vccd1 _4705_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5138__A _5975_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4636_ _5692_/Q _5669_/Q _4645_/S vssd1 vssd1 vccd1 vccd1 _4636_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4567_ _4567_/A vssd1 vssd1 vccd1 vccd1 _4567_/Y sky130_fd_sc_hd__inv_2
X_4498_ _3561_/A _3542_/A _5864_/Q vssd1 vssd1 vccd1 vccd1 _4502_/B sky130_fd_sc_hd__a21oi_1
X_3518_ _3518_/A _3518_/B vssd1 vssd1 vccd1 vccd1 _3518_/Y sky130_fd_sc_hd__nor2_1
XFILLER_1_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3449_ _3896_/A _3469_/B _2928_/B _3448_/Y vssd1 vssd1 vccd1 vccd1 _3449_/X sky130_fd_sc_hd__a2bb2o_1
XANTENNA__4188__S _4200_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5119_ _5069_/X _5104_/A _5118_/X _5114_/X vssd1 vssd1 vccd1 vccd1 _5968_/D sky130_fd_sc_hd__o211a_1
XFILLER_17_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6099_ _6101_/CLK _6099_/D vssd1 vssd1 vccd1 vccd1 _6099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2960__A _3518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3031__A _3897_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3966__A _3966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5470_ _5470_/A vssd1 vssd1 vccd1 vccd1 _5470_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5173__C1 _5172_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4421_ _5842_/Q _4419_/X _4433_/S vssd1 vssd1 vccd1 vccd1 _4422_/A sky130_fd_sc_hd__mux2_1
X_4352_ _4352_/A vssd1 vssd1 vccd1 vccd1 _5821_/D sky130_fd_sc_hd__clkbuf_1
X_3303_ _3428_/A vssd1 vssd1 vccd1 vccd1 _3486_/A sky130_fd_sc_hd__clkbuf_2
X_4283_ _4283_/A _4283_/B _4283_/C vssd1 vssd1 vccd1 vccd1 _4283_/X sky130_fd_sc_hd__or3_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5405__B _5405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3206__A _6020_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3234_ _6031_/Q _5932_/Q vssd1 vssd1 vccd1 vccd1 _3234_/Y sky130_fd_sc_hd__xnor2_1
X_6022_ _6024_/CLK _6022_/D vssd1 vssd1 vccd1 vccd1 _6022_/Q sky130_fd_sc_hd__dfxtp_1
Xuser_proj_example_99 vssd1 vssd1 vccd1 vccd1 user_proj_example_99/HI io_oeb[17] sky130_fd_sc_hd__conb_1
Xuser_proj_example_88 vssd1 vssd1 vccd1 vccd1 user_proj_example_88/HI io_oeb[6] sky130_fd_sc_hd__conb_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3165_ _3079_/B _3350_/C _3341_/B _3071_/A vssd1 vssd1 vccd1 vccd1 _3165_/X sky130_fd_sc_hd__a22o_1
X_3096_ _3928_/A vssd1 vssd1 vccd1 vccd1 _3814_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5806_ _5808_/CLK _5806_/D vssd1 vssd1 vccd1 vccd1 _5806_/Q sky130_fd_sc_hd__dfxtp_1
X_3998_ _3938_/A _3932_/A _3997_/X vssd1 vssd1 vccd1 vccd1 _3999_/B sky130_fd_sc_hd__a21oi_1
XFILLER_10_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5737_ _6121_/CLK _5737_/D vssd1 vssd1 vccd1 vccd1 _5737_/Q sky130_fd_sc_hd__dfxtp_1
X_2949_ _3312_/C _3312_/D _2949_/C _2949_/D vssd1 vssd1 vccd1 vccd1 _3296_/B sky130_fd_sc_hd__or4_4
XFILLER_13_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5668_ _6091_/CLK _5668_/D vssd1 vssd1 vccd1 vccd1 _5668_/Q sky130_fd_sc_hd__dfxtp_1
X_4619_ _5126_/A vssd1 vssd1 vccd1 vccd1 _4824_/A sky130_fd_sc_hd__clkbuf_2
X_5599_ _6104_/Q _5599_/B vssd1 vssd1 vccd1 vccd1 _5599_/X sky130_fd_sc_hd__or2_1
XFILLER_89_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2955__A _3296_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3786__A _4251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_531 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3001__D _3440_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_1_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6048_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__2849__B _5736_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_43_wb_clk_i_A clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_5_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output57_A _5884_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4970_ _4970_/A _4970_/B _4970_/C vssd1 vssd1 vccd1 vccd1 _4971_/A sky130_fd_sc_hd__and3_1
XFILLER_63_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3921_ _4010_/A _3921_/B _3921_/C vssd1 vssd1 vccd1 vccd1 _3922_/S sky130_fd_sc_hd__and3b_1
XFILLER_44_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3852_ _5241_/B _4218_/A vssd1 vssd1 vccd1 vccd1 _3897_/D sky130_fd_sc_hd__nand2_1
X_3783_ _3611_/A _5710_/Q _3791_/S vssd1 vssd1 vccd1 vccd1 _3784_/B sky130_fd_sc_hd__mux2_1
X_5522_ _6075_/Q _5526_/B vssd1 vssd1 vccd1 vccd1 _5522_/X sky130_fd_sc_hd__or2_1
X_5453_ _5376_/X _5449_/X _5452_/X _5446_/X vssd1 vssd1 vccd1 vccd1 _6049_/D sky130_fd_sc_hd__o211a_1
X_4404_ _4402_/A _5254_/C _5837_/Q vssd1 vssd1 vccd1 vccd1 _4404_/X sky130_fd_sc_hd__o21a_1
X_5384_ _5384_/A _5387_/B vssd1 vssd1 vccd1 vccd1 _5384_/Y sky130_fd_sc_hd__nand2_1
X_4335_ _3322_/X _4337_/S _4333_/Y _6066_/Q vssd1 vssd1 vccd1 vccd1 _5815_/D sky130_fd_sc_hd__a22o_1
XFILLER_59_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4266_ _4321_/S _3480_/C _4294_/A vssd1 vssd1 vccd1 vccd1 _4269_/B sky130_fd_sc_hd__o21ba_1
X_3217_ _4954_/A vssd1 vssd1 vccd1 vccd1 _4972_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6005_ _6005_/CLK _6005_/D vssd1 vssd1 vccd1 vccd1 _6005_/Q sky130_fd_sc_hd__dfxtp_1
X_4197_ _5801_/Q _4196_/X _4200_/S vssd1 vssd1 vccd1 vccd1 _4198_/A sky130_fd_sc_hd__mux2_1
X_3148_ _5988_/Q vssd1 vssd1 vccd1 vccd1 _4480_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_39_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3079_ _3266_/A _3079_/B vssd1 vssd1 vccd1 vccd1 _3079_/X sky130_fd_sc_hd__and2_1
XFILLER_54_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_87 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4663__A1 _5882_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4120_ _5778_/Q _4118_/X _4133_/S vssd1 vssd1 vccd1 vccd1 _4121_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4051_ _4051_/A vssd1 vssd1 vccd1 vccd1 _5758_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3002_ _3476_/C _2973_/X _2984_/X _2991_/X _3001_/X vssd1 vssd1 vccd1 vccd1 _3022_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_49_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput5 la_data_in[32] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4953_ _4953_/A _4953_/B vssd1 vssd1 vccd1 vccd1 _4958_/B sky130_fd_sc_hd__nor2_1
XFILLER_17_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3904_ _3895_/X _3287_/X _3904_/S vssd1 vssd1 vccd1 vccd1 _3905_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4884_ _5958_/Q _4882_/X _4916_/S vssd1 vssd1 vccd1 vccd1 _4884_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3835_ _4218_/A _3283_/B _3553_/A vssd1 vssd1 vccd1 vccd1 _4288_/A sky130_fd_sc_hd__a21o_1
X_3766_ _3791_/S vssd1 vssd1 vccd1 vccd1 _3780_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__4590__A0 _6113_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5505_ _6069_/Q _5505_/B vssd1 vssd1 vccd1 vccd1 _5505_/X sky130_fd_sc_hd__or2_1
X_3697_ _3607_/A _5686_/Q _3697_/S vssd1 vssd1 vccd1 vccd1 _3698_/B sky130_fd_sc_hd__mux2_1
XFILLER_10_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5436_ _5357_/X _5427_/X _5434_/X _5435_/X vssd1 vssd1 vccd1 vccd1 _6043_/D sky130_fd_sc_hd__o211a_1
XFILLER_87_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5367_ _6022_/Q _5367_/B vssd1 vssd1 vccd1 vccd1 _5367_/X sky130_fd_sc_hd__or2_1
X_5298_ _5297_/A _5323_/A vssd1 vssd1 vccd1 vccd1 _5299_/B sky130_fd_sc_hd__and2b_1
X_4318_ _5301_/C _3880_/X _4317_/X _3111_/X vssd1 vssd1 vccd1 vccd1 _4318_/X sky130_fd_sc_hd__a211o_1
X_4249_ _5806_/Q _4249_/B _4249_/C vssd1 vssd1 vccd1 vccd1 _4275_/C sky130_fd_sc_hd__and3_1
XFILLER_74_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3384__B2 _4366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5056__A _5056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5530__C1 _5529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3304__A _3480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3620_ _5046_/A _5046_/B _3620_/C vssd1 vssd1 vccd1 vccd1 _5343_/B sky130_fd_sc_hd__and3_2
X_3551_ _5667_/Q _5713_/Q _4562_/B vssd1 vssd1 vccd1 vccd1 _3551_/X sky130_fd_sc_hd__and3b_1
X_3482_ _3482_/A _3482_/B vssd1 vssd1 vccd1 vccd1 _3482_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5221_ _5221_/A vssd1 vssd1 vccd1 vccd1 _6002_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5152_ _5979_/Q _5162_/B vssd1 vssd1 vccd1 vccd1 _5152_/X sky130_fd_sc_hd__or2_1
X_4103_ _4103_/A vssd1 vssd1 vccd1 vccd1 _5773_/D sky130_fd_sc_hd__clkbuf_1
X_5083_ _5955_/Q _5093_/B vssd1 vssd1 vccd1 vccd1 _5083_/X sky130_fd_sc_hd__or2_1
X_4034_ _4034_/A vssd1 vssd1 vccd1 vccd1 _5753_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5985_ _6003_/CLK _5985_/D vssd1 vssd1 vccd1 vccd1 _5985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4936_ _6039_/Q _4924_/X _4935_/Y _4929_/X vssd1 vssd1 vccd1 vccd1 _5913_/D sky130_fd_sc_hd__o211a_1
X_4867_ _5980_/Q _4854_/X _4855_/X vssd1 vssd1 vccd1 vccd1 _4867_/X sky130_fd_sc_hd__o21a_1
XFILLER_20_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3818_ _5337_/S _5716_/Q vssd1 vssd1 vccd1 vccd1 _3818_/X sky130_fd_sc_hd__and2b_1
X_4798_ _5661_/Q _4797_/X _4821_/S vssd1 vssd1 vccd1 vccd1 _4798_/X sky130_fd_sc_hd__mux2_1
X_3749_ _5389_/A _5700_/Q _3753_/S vssd1 vssd1 vccd1 vccd1 _3750_/B sky130_fd_sc_hd__mux2_1
XFILLER_4_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5419_ _6038_/Q _5424_/B vssd1 vssd1 vccd1 vccd1 _5419_/X sky130_fd_sc_hd__or2_1
XFILLER_47_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_proj_example_103 vssd1 vssd1 vccd1 vccd1 user_proj_example_103/HI io_oeb[21]
+ sky130_fd_sc_hd__conb_1
XANTENNA__3794__A _3794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_proj_example_114 vssd1 vssd1 vccd1 vccd1 user_proj_example_114/HI io_oeb[32]
+ sky130_fd_sc_hd__conb_1
XANTENNA__4554__A0 _5665_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xuser_proj_example_125 vssd1 vssd1 vccd1 vccd1 user_proj_example_125/HI la_data_out[0]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_136 vssd1 vssd1 vccd1 vccd1 user_proj_example_136/HI la_data_out[11]
+ sky130_fd_sc_hd__conb_1
XANTENNA__4402__B _5254_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xuser_proj_example_169 vssd1 vssd1 vccd1 vccd1 user_proj_example_169/HI la_data_out[44]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_147 vssd1 vssd1 vccd1 vccd1 user_proj_example_147/HI la_data_out[22]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_158 vssd1 vssd1 vccd1 vccd1 user_proj_example_158/HI la_data_out[33]
+ sky130_fd_sc_hd__conb_1
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4609__A1 _5877_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2982_ _4218_/B _2982_/B vssd1 vssd1 vccd1 vccd1 _2983_/B sky130_fd_sc_hd__nand2_1
X_5770_ _5914_/CLK _5770_/D vssd1 vssd1 vccd1 vccd1 _5770_/Q sky130_fd_sc_hd__dfxtp_1
X_4721_ _6076_/Q _4732_/B vssd1 vssd1 vccd1 vccd1 _4721_/X sky130_fd_sc_hd__or2_1
X_4652_ _5881_/Q _4579_/X _4650_/X _4651_/X vssd1 vssd1 vccd1 vccd1 _5881_/D sky130_fd_sc_hd__a22o_1
Xinput30 la_data_in[55] vssd1 vssd1 vccd1 vccd1 _3617_/A sky130_fd_sc_hd__clkbuf_1
X_3603_ _3601_/X _3592_/X _3602_/X _3585_/X vssd1 vssd1 vccd1 vccd1 _5660_/D sky130_fd_sc_hd__o211a_1
Xinput41 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 _3570_/B sky130_fd_sc_hd__clkbuf_1
X_4583_ _4859_/A vssd1 vssd1 vccd1 vccd1 _4706_/A sky130_fd_sc_hd__clkbuf_2
X_3534_ _5868_/Q vssd1 vssd1 vccd1 vccd1 _4545_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3465_ _2959_/C _3465_/B _3465_/C vssd1 vssd1 vccd1 vccd1 _3840_/B sky130_fd_sc_hd__nand3b_1
X_5204_ _5204_/A _5204_/B vssd1 vssd1 vccd1 vccd1 _5205_/A sky130_fd_sc_hd__and2_1
XANTENNA__5424__A _6040_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3396_ _5234_/A _4293_/A vssd1 vssd1 vccd1 vccd1 _3396_/Y sky130_fd_sc_hd__nor2_1
XFILLER_69_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5135_ _5059_/X _5125_/X _5134_/X _5130_/X vssd1 vssd1 vccd1 vccd1 _5973_/D sky130_fd_sc_hd__o211a_1
XFILLER_29_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5066_ _5951_/Q _5066_/B vssd1 vssd1 vccd1 vccd1 _5066_/X sky130_fd_sc_hd__or2_1
XANTENNA__5273__A1 _5301_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4017_ _4017_/A vssd1 vssd1 vccd1 vccd1 _4017_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5968_ _5975_/CLK _5968_/D vssd1 vssd1 vccd1 vccd1 _5968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_404 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4919_ _5978_/Q _4706_/A _4716_/A _4918_/X vssd1 vssd1 vccd1 vccd1 _4919_/X sky130_fd_sc_hd__a211o_1
X_5899_ _6088_/CLK _5899_/D vssd1 vssd1 vccd1 vccd1 _5899_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3511__A1 _3269_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4384__S _4396_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input19_A la_data_in[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3789__A _3966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3029__A _3826_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2868__A _3459_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ _3247_/Y _5852_/Q _5171_/A vssd1 vssd1 vccd1 vccd1 _5852_/D sky130_fd_sc_hd__a21o_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3181_ _5925_/Q vssd1 vssd1 vccd1 vccd1 _3186_/A sky130_fd_sc_hd__inv_2
XFILLER_66_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5822_ _6048_/CLK _5822_/D vssd1 vssd1 vccd1 vccd1 _5822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5753_ _5796_/CLK _5753_/D vssd1 vssd1 vccd1 vccd1 _5753_/Q sky130_fd_sc_hd__dfxtp_1
X_2965_ _3850_/C _2972_/C vssd1 vssd1 vccd1 vccd1 _4229_/A sky130_fd_sc_hd__or2_2
X_4704_ _5886_/Q _4653_/X _4702_/X _4703_/Y vssd1 vssd1 vccd1 vccd1 _5886_/D sky130_fd_sc_hd__a22o_1
XANTENNA__5419__A _6038_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2896_ _2896_/A vssd1 vssd1 vccd1 vccd1 _5279_/A sky130_fd_sc_hd__clkbuf_2
X_5684_ _6085_/CLK _5684_/D vssd1 vssd1 vccd1 vccd1 _5684_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4635_ _5879_/Q _4579_/X _4633_/X _4634_/X vssd1 vssd1 vccd1 vccd1 _5879_/D sky130_fd_sc_hd__a22o_1
X_4566_ _5188_/A vssd1 vssd1 vccd1 vccd1 _5186_/A sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_25_wb_clk_i clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5945_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3517_ _3374_/A _3513_/B _3071_/A vssd1 vssd1 vccd1 vccd1 _3517_/X sky130_fd_sc_hd__a21o_1
X_4497_ _4496_/Y _5857_/Q _3529_/B _4568_/B vssd1 vssd1 vccd1 vccd1 _4502_/A sky130_fd_sc_hd__o31a_1
XANTENNA__5154__A _5980_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3448_ _3448_/A vssd1 vssd1 vccd1 vccd1 _3448_/Y sky130_fd_sc_hd__clkinv_2
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3379_ _3379_/A vssd1 vssd1 vccd1 vccd1 _4450_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_57_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5118_ _5968_/Q _5122_/B vssd1 vssd1 vccd1 vccd1 _5118_/X sky130_fd_sc_hd__or2_1
X_6098_ _6138_/CLK _6098_/D vssd1 vssd1 vccd1 vccd1 _6098_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5601__B _5601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5049_ _5622_/A _5148_/B vssd1 vssd1 vccd1 vccd1 _5050_/A sky130_fd_sc_hd__or2_1
XFILLER_72_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2960__B _3283_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_278 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5182__A0 _5059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_33_wb_clk_i_A clkbuf_3_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_4_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5237__A1 _3480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_123 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4212__A2 _3839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4420_ _4420_/A vssd1 vssd1 vccd1 vccd1 _4433_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_8_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4920__B1 _4607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4351_ _5821_/Q _4350_/X _4357_/S vssd1 vssd1 vccd1 vccd1 _4352_/A sky130_fd_sc_hd__mux2_1
X_3302_ _4255_/A vssd1 vssd1 vccd1 vccd1 _3428_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4282_ _5247_/A _3282_/A _3850_/C _4281_/D _4471_/B vssd1 vssd1 vccd1 vccd1 _4282_/X
+ sky130_fd_sc_hd__o41a_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3233_ _6029_/Q _5930_/Q vssd1 vssd1 vccd1 vccd1 _3233_/X sky130_fd_sc_hd__and2_1
X_6021_ _6024_/CLK _6021_/D vssd1 vssd1 vccd1 vccd1 _6021_/Q sky130_fd_sc_hd__dfxtp_1
Xuser_proj_example_89 vssd1 vssd1 vccd1 vccd1 user_proj_example_89/HI io_oeb[7] sky130_fd_sc_hd__conb_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3164_ _3839_/A _4321_/S vssd1 vssd1 vccd1 vccd1 _3341_/B sky130_fd_sc_hd__nor2_1
X_3095_ _3838_/A vssd1 vssd1 vccd1 vccd1 _3928_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_81_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4739__A0 _6102_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5805_ _5808_/CLK _5805_/D vssd1 vssd1 vccd1 vccd1 _5805_/Q sky130_fd_sc_hd__dfxtp_1
X_3997_ _5735_/Q _3941_/A _3945_/X _3996_/Y vssd1 vssd1 vccd1 vccd1 _3997_/X sky130_fd_sc_hd__o211a_1
XANTENNA__5400__A1 _3563_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2948_ _3849_/B _3003_/A _5247_/B _3434_/A vssd1 vssd1 vccd1 vccd1 _2948_/X sky130_fd_sc_hd__a22o_1
X_5736_ _5736_/CLK _5736_/D vssd1 vssd1 vccd1 vccd1 _5736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5667_ _6024_/CLK _5667_/D vssd1 vssd1 vccd1 vccd1 _5667_/Q sky130_fd_sc_hd__dfxtp_2
X_2879_ _5813_/Q vssd1 vssd1 vccd1 vccd1 _3838_/A sky130_fd_sc_hd__clkbuf_2
X_4618_ _6066_/Q _5537_/B vssd1 vssd1 vccd1 vccd1 _4618_/X sky130_fd_sc_hd__or2_1
X_5598_ _3563_/X _5580_/A _5596_/X _5597_/X vssd1 vssd1 vccd1 vccd1 _6103_/D sky130_fd_sc_hd__o211a_1
X_4549_ _4549_/A _4549_/B vssd1 vssd1 vccd1 vccd1 _5870_/D sky130_fd_sc_hd__nor2_1
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4199__S _4554_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5612__A _5638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2955__B _5327_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5059__A _5059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3920_ _6120_/Q _3491_/X _3919_/X vssd1 vssd1 vccd1 vccd1 _3920_/X sky130_fd_sc_hd__o21a_1
XFILLER_51_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5630__A1 _5353_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3641__A0 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3851_ _5250_/A _4470_/C _3851_/C _3851_/D vssd1 vssd1 vccd1 vccd1 _3913_/B sky130_fd_sc_hd__and4_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3782_ _3782_/A vssd1 vssd1 vccd1 vccd1 _5709_/D sky130_fd_sc_hd__clkbuf_1
X_5521_ _5382_/X _5514_/X _5520_/X _5518_/X vssd1 vssd1 vccd1 vccd1 _6074_/D sky130_fd_sc_hd__o211a_1
X_5452_ _6049_/Q _5460_/B vssd1 vssd1 vccd1 vccd1 _5452_/X sky130_fd_sc_hd__or2_1
X_4403_ _4420_/A vssd1 vssd1 vccd1 vccd1 _4417_/S sky130_fd_sc_hd__clkbuf_2
X_5383_ _5401_/B vssd1 vssd1 vccd1 vccd1 _5387_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4334_ _3438_/A _4337_/S _4333_/Y _6065_/Q vssd1 vssd1 vccd1 vccd1 _5814_/D sky130_fd_sc_hd__a22o_1
XFILLER_5_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4265_ _4233_/A _3266_/Y _4264_/X vssd1 vssd1 vccd1 vccd1 _4270_/B sky130_fd_sc_hd__o21ai_1
X_6004_ _6087_/CLK _6004_/D vssd1 vssd1 vccd1 vccd1 _6004_/Q sky130_fd_sc_hd__dfxtp_1
X_3216_ _5873_/Q _5852_/Q vssd1 vssd1 vccd1 vccd1 _4942_/B sky130_fd_sc_hd__and2_1
XFILLER_39_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4196_ _5951_/Q _5800_/Q _4196_/S vssd1 vssd1 vccd1 vccd1 _4196_/X sky130_fd_sc_hd__mux2_1
X_3147_ _4567_/A _3147_/B vssd1 vssd1 vccd1 vccd1 _3546_/A sky130_fd_sc_hd__or2_1
XFILLER_67_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3078_ _5255_/A vssd1 vssd1 vccd1 vccd1 _3079_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_35_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_40_wb_clk_i clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5966_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_5719_ _6067_/CLK _5719_/D vssd1 vssd1 vccd1 vccd1 _5719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5342__A input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3797__A _4855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3926__A1 _4210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3037__A _3037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4050_ _5758_/Q _4048_/X _4063_/S vssd1 vssd1 vccd1 vccd1 _4051_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3001_ _3484_/A _5301_/B _3440_/B _3440_/C vssd1 vssd1 vccd1 vccd1 _3001_/X sky130_fd_sc_hd__and4bb_1
XANTENNA__3457__A3 _3326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_462 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput6 la_data_in[33] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5064__C1 _5043_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4952_ _4953_/A _4953_/B vssd1 vssd1 vccd1 vccd1 _4957_/A sky130_fd_sc_hd__and2_1
X_3903_ _3903_/A _3913_/A _3903_/C _5261_/B vssd1 vssd1 vccd1 vccd1 _3904_/S sky130_fd_sc_hd__or4_1
X_4883_ _4883_/A vssd1 vssd1 vccd1 vccd1 _4916_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_32_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3834_ _3834_/A _3834_/B vssd1 vssd1 vccd1 vccd1 _5254_/A sky130_fd_sc_hd__and2_1
XFILLER_32_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3765_ _3765_/A _5201_/A vssd1 vssd1 vccd1 vccd1 _3791_/S sky130_fd_sc_hd__nand2_1
XANTENNA__3873__C _3873_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3696_ _3696_/A vssd1 vssd1 vccd1 vccd1 _5685_/D sky130_fd_sc_hd__clkbuf_1
X_5504_ _5360_/X _5493_/X _5502_/X _5503_/X vssd1 vssd1 vccd1 vccd1 _6068_/D sky130_fd_sc_hd__o211a_1
X_5435_ _5461_/A vssd1 vssd1 vccd1 vccd1 _5435_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4342__A1 _4366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5366_ _5366_/A vssd1 vssd1 vccd1 vccd1 _5366_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_87_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5297_ _5297_/A _5297_/B _5297_/C vssd1 vssd1 vccd1 vccd1 _5310_/A sky130_fd_sc_hd__and3_1
X_4317_ _3494_/B _5304_/B _3869_/X _3867_/X vssd1 vssd1 vccd1 vccd1 _4317_/X sky130_fd_sc_hd__o211a_1
X_4248_ _4249_/B _4228_/X _5806_/Q vssd1 vssd1 vccd1 vccd1 _4250_/B sky130_fd_sc_hd__a21oi_1
XFILLER_74_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4179_ _5664_/Q _5795_/Q _4179_/S vssd1 vssd1 vccd1 vccd1 _4179_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5055__C1 _5043_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4387__S _4396_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3550_ _5945_/Q _5741_/Q vssd1 vssd1 vccd1 vccd1 _3550_/X sky130_fd_sc_hd__and2b_1
X_3481_ _4438_/A _3481_/B vssd1 vssd1 vccd1 vccd1 _3482_/B sky130_fd_sc_hd__or2_1
X_5220_ _5220_/A _5220_/B vssd1 vssd1 vccd1 vccd1 _5221_/A sky130_fd_sc_hd__and2_1
XFILLER_69_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5151_ _5168_/B vssd1 vssd1 vccd1 vccd1 _5162_/B sky130_fd_sc_hd__clkbuf_1
X_4102_ _5773_/Q _4099_/X _4116_/S vssd1 vssd1 vccd1 vccd1 _4103_/A sky130_fd_sc_hd__mux2_1
X_5082_ _5100_/B vssd1 vssd1 vccd1 vccd1 _5093_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_84_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4033_ _5753_/Q _4030_/X _4046_/S vssd1 vssd1 vccd1 vccd1 _4034_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3835__B1 _3553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5984_ _6003_/CLK _5984_/D vssd1 vssd1 vccd1 vccd1 _5984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3230__A _6033_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4935_ _4935_/A _4944_/B vssd1 vssd1 vccd1 vccd1 _4935_/Y sky130_fd_sc_hd__nand2_1
X_4866_ _5972_/Q _4859_/X _4818_/X _4865_/X vssd1 vssd1 vccd1 vccd1 _4866_/X sky130_fd_sc_hd__a211o_1
X_3817_ _5340_/S vssd1 vssd1 vccd1 vccd1 _5337_/S sky130_fd_sc_hd__dlymetal6s2s_1
X_4797_ _5708_/Q _5685_/Q _4797_/S vssd1 vssd1 vccd1 vccd1 _4797_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4061__A _4095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3748_ _3748_/A vssd1 vssd1 vccd1 vccd1 _5699_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5157__A _5408_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3679_ _3684_/A _3679_/B vssd1 vssd1 vccd1 vccd1 _3680_/A sky130_fd_sc_hd__and2_1
X_5418_ _3607_/X _5404_/X _5417_/X _5409_/X vssd1 vssd1 vccd1 vccd1 _6037_/D sky130_fd_sc_hd__o211a_1
X_5349_ _5405_/B _5622_/B vssd1 vssd1 vccd1 vccd1 _5374_/B sky130_fd_sc_hd__nor2_1
XFILLER_87_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5620__A _6112_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3140__A _3411_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xuser_proj_example_115 vssd1 vssd1 vccd1 vccd1 user_proj_example_115/HI io_oeb[33]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_104 vssd1 vssd1 vccd1 vccd1 user_proj_example_104/HI io_oeb[22]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_126 vssd1 vssd1 vccd1 vccd1 user_proj_example_126/HI la_data_out[1]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_137 vssd1 vssd1 vccd1 vccd1 user_proj_example_137/HI la_data_out[12]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_159 vssd1 vssd1 vccd1 vccd1 user_proj_example_159/HI la_data_out[34]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_148 vssd1 vssd1 vccd1 vccd1 user_proj_example_148/HI la_data_out[23]
+ sky130_fd_sc_hd__conb_1
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5813__CLK _5813_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2981_ _3824_/A _5718_/Q vssd1 vssd1 vccd1 vccd1 _2982_/B sky130_fd_sc_hd__xor2_2
XFILLER_21_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4720_ _6100_/Q _4719_/X _4720_/S vssd1 vssd1 vccd1 vccd1 _4720_/X sky130_fd_sc_hd__mux2_1
XFILLER_42_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4651_ _6021_/Q _4606_/X _4607_/X vssd1 vssd1 vccd1 vccd1 _4651_/X sky130_fd_sc_hd__o21a_1
Xinput20 la_data_in[46] vssd1 vssd1 vccd1 vccd1 _3563_/A sky130_fd_sc_hd__clkbuf_1
Xinput31 la_data_in[56] vssd1 vssd1 vccd1 vccd1 _5045_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3602_ _5660_/Q _3608_/B vssd1 vssd1 vccd1 vccd1 _3602_/X sky130_fd_sc_hd__or2_1
Xinput42 wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 _3564_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4582_ _4597_/A _4604_/B vssd1 vssd1 vccd1 vccd1 _4859_/A sky130_fd_sc_hd__nor2_2
X_3533_ _5859_/Q _5858_/Q _3147_/B vssd1 vssd1 vccd1 vccd1 _3544_/B sky130_fd_sc_hd__o21bai_1
XFILLER_6_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3464_ _3837_/A _3040_/B _3463_/X vssd1 vssd1 vccd1 vccd1 _3464_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_88_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5203_ _5045_/A _5997_/Q _5216_/S vssd1 vssd1 vccd1 vccd1 _5204_/B sky130_fd_sc_hd__mux2_1
X_3395_ _5714_/Q _3826_/C vssd1 vssd1 vccd1 vccd1 _3800_/B sky130_fd_sc_hd__nor2_1
X_5134_ _5973_/Q _5138_/B vssd1 vssd1 vccd1 vccd1 _5134_/X sky130_fd_sc_hd__or2_1
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5065_ _5065_/A vssd1 vssd1 vccd1 vccd1 _5065_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3284__A1 _3117_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4016_ _4113_/A _4016_/B vssd1 vssd1 vccd1 vccd1 _4017_/A sky130_fd_sc_hd__and2_1
XFILLER_25_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5967_ _5975_/CLK _5967_/D vssd1 vssd1 vccd1 vccd1 _5967_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4918_ _4717_/A _4916_/X _4917_/X _5469_/B vssd1 vssd1 vccd1 vccd1 _4918_/X sky130_fd_sc_hd__o211a_1
XFILLER_33_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5898_ _6088_/CLK _5898_/D vssd1 vssd1 vccd1 vccd1 _5898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4849_ _5947_/Q _4848_/X _4872_/S vssd1 vssd1 vccd1 vccd1 _4849_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_23_wb_clk_i_A clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__5497__C1 _5488_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3135__A _3135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5836__CLK _5836_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5421__C1 _5420_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3045__A _3857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3180_ _5926_/Q vssd1 vssd1 vccd1 vccd1 _3180_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5821_ _6117_/CLK _5821_/D vssd1 vssd1 vccd1 vccd1 _5821_/Q sky130_fd_sc_hd__dfxtp_1
X_2964_ _3038_/A _5717_/Q vssd1 vssd1 vccd1 vccd1 _2972_/C sky130_fd_sc_hd__xor2_1
X_5752_ _5796_/CLK _5752_/D vssd1 vssd1 vccd1 vccd1 _5752_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4703_ _5384_/A _4602_/X _4623_/X vssd1 vssd1 vccd1 vccd1 _4703_/Y sky130_fd_sc_hd__a21oi_1
X_2895_ _5872_/Q vssd1 vssd1 vccd1 vccd1 _2896_/A sky130_fd_sc_hd__inv_2
X_5683_ _6085_/CLK _5683_/D vssd1 vssd1 vccd1 vccd1 _5683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4634_ _6019_/Q _4606_/X _4607_/X vssd1 vssd1 vccd1 vccd1 _4634_/X sky130_fd_sc_hd__o21a_1
X_4565_ _3135_/A _5743_/Q _4562_/X _4564_/X vssd1 vssd1 vccd1 vccd1 _5874_/D sky130_fd_sc_hd__a31o_1
X_3516_ _2899_/A _3291_/B _3513_/B _3410_/X vssd1 vssd1 vccd1 vccd1 _3516_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5435__A _5461_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4496_ _5988_/Q vssd1 vssd1 vccd1 vccd1 _4496_/Y sky130_fd_sc_hd__inv_2
X_3447_ _3857_/B _3047_/X _2936_/A _3880_/S vssd1 vssd1 vccd1 vccd1 _3447_/X sky130_fd_sc_hd__a22o_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3378_ _6121_/Q vssd1 vssd1 vccd1 vccd1 _3379_/A sky130_fd_sc_hd__clkbuf_2
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6097_ _6135_/CLK _6097_/D vssd1 vssd1 vccd1 vccd1 _6097_/Q sky130_fd_sc_hd__dfxtp_1
X_5117_ _5065_/X _5104_/X _5116_/X _5114_/X vssd1 vssd1 vccd1 vccd1 _5967_/D sky130_fd_sc_hd__o211a_1
XFILLER_84_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5048_ _5051_/A vssd1 vssd1 vccd1 vccd1 _5148_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_27_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5651__C1 _5172_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4233__B _4233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input31_A la_data_in[56] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5255__A _5255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4350_ _6043_/Q _5820_/Q _4363_/S vssd1 vssd1 vccd1 vccd1 _4350_/X sky130_fd_sc_hd__mux2_1
X_3301_ _4458_/A _3284_/Y _3291_/X _3300_/X vssd1 vssd1 vccd1 vccd1 _3301_/X sky130_fd_sc_hd__a211o_1
X_4281_ _4281_/A _5720_/Q _4281_/C _4281_/D vssd1 vssd1 vccd1 vccd1 _4471_/B sky130_fd_sc_hd__or4_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3232_ _6029_/Q _5930_/Q vssd1 vssd1 vccd1 vccd1 _3232_/Y sky130_fd_sc_hd__nor2_1
X_6020_ _6024_/CLK _6020_/D vssd1 vssd1 vccd1 vccd1 _6020_/Q sky130_fd_sc_hd__dfxtp_1
X_3163_ _5836_/Q vssd1 vssd1 vccd1 vccd1 _4321_/S sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3094_ _3391_/A vssd1 vssd1 vccd1 vccd1 _3135_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_54_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3239__A1 _5401_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3239__B2 _5384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5804_ _6131_/CLK _5804_/D vssd1 vssd1 vccd1 vccd1 _5804_/Q sky130_fd_sc_hd__dfxtp_1
X_3996_ _5735_/Q _3996_/B vssd1 vssd1 vccd1 vccd1 _3996_/Y sky130_fd_sc_hd__nand2_1
XFILLER_22_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2947_ _5285_/A _3400_/B vssd1 vssd1 vccd1 vccd1 _3434_/A sky130_fd_sc_hd__nor2_2
X_5735_ _5808_/CLK _5735_/D vssd1 vssd1 vccd1 vccd1 _5735_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5666_ _6018_/CLK _5666_/D vssd1 vssd1 vccd1 vccd1 _5666_/Q sky130_fd_sc_hd__dfxtp_2
X_2878_ _2944_/B _4464_/B vssd1 vssd1 vccd1 vccd1 _3833_/C sky130_fd_sc_hd__or2_1
X_4617_ _5102_/A vssd1 vssd1 vccd1 vccd1 _5537_/B sky130_fd_sc_hd__clkbuf_2
X_5597_ _5597_/A vssd1 vssd1 vccd1 vccd1 _5597_/X sky130_fd_sc_hd__clkbuf_2
X_4548_ _4548_/A _4548_/B vssd1 vssd1 vccd1 vccd1 _4549_/B sky130_fd_sc_hd__xnor2_1
X_4479_ _3336_/X _4281_/D _4478_/X vssd1 vssd1 vccd1 vccd1 _5856_/D sky130_fd_sc_hd__o21a_1
XFILLER_1_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2955__C _2955_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3307__B _3857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2881__B _3836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3850_ _4470_/A _4470_/B _3850_/C vssd1 vssd1 vccd1 vccd1 _3851_/D sky130_fd_sc_hd__and3_1
X_3781_ _3784_/A _3781_/B vssd1 vssd1 vccd1 vccd1 _3782_/A sky130_fd_sc_hd__and2_1
X_5520_ _6074_/Q _5526_/B vssd1 vssd1 vccd1 vccd1 _5520_/X sky130_fd_sc_hd__or2_1
XFILLER_8_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5451_ _5467_/B vssd1 vssd1 vccd1 vccd1 _5460_/B sky130_fd_sc_hd__clkbuf_1
X_4402_ _4402_/A _5254_/C vssd1 vssd1 vccd1 vccd1 _4420_/A sky130_fd_sc_hd__nor2_1
X_5382_ _5382_/A vssd1 vssd1 vccd1 vccd1 _5382_/X sky130_fd_sc_hd__buf_2
X_4333_ _6068_/Q _4337_/S vssd1 vssd1 vccd1 vccd1 _4333_/Y sky130_fd_sc_hd__nor2_1
XFILLER_5_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4264_ _3276_/Y _4294_/B _4242_/C _3800_/B vssd1 vssd1 vccd1 vccd1 _4264_/X sky130_fd_sc_hd__o22a_1
X_3215_ _4946_/C _4954_/A _3215_/C vssd1 vssd1 vccd1 vccd1 _5011_/B sky130_fd_sc_hd__and3_1
X_6003_ _6003_/CLK _6003_/D vssd1 vssd1 vccd1 vccd1 _6003_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4657__A0 _6118_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4195_ _4195_/A vssd1 vssd1 vccd1 vccd1 _5800_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3233__A _6029_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3146_ _5850_/Q _3146_/B vssd1 vssd1 vccd1 vccd1 _3147_/B sky130_fd_sc_hd__xnor2_1
XFILLER_82_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3077_ _3824_/D vssd1 vssd1 vccd1 vccd1 _5255_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_54_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5606__C1 _5597_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5385__A1 _5382_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3979_ _3979_/A _3979_/B vssd1 vssd1 vccd1 vccd1 _5730_/D sky130_fd_sc_hd__nor2_1
X_5718_ _5796_/CLK _5718_/D vssd1 vssd1 vccd1 vccd1 _5718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5649_ _5386_/X _3576_/X _5648_/X _5172_/X vssd1 vssd1 vccd1 vccd1 _6135_/D sky130_fd_sc_hd__o211a_1
XFILLER_40_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_1__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2982__A _4218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3871__A1 _3873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output62_A _5889_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3000_ _3297_/B _3891_/A vssd1 vssd1 vccd1 vccd1 _3440_/C sky130_fd_sc_hd__nor2_1
XFILLER_64_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput7 la_data_in[34] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2892__A _3480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3862__A1 _3484_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4951_ _5918_/Q _4948_/X _4953_/B _4940_/X vssd1 vssd1 vccd1 vccd1 _5918_/D sky130_fd_sc_hd__o211a_1
XFILLER_24_319 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3902_ _5233_/B _3902_/B _3902_/C _3901_/Y vssd1 vssd1 vccd1 vccd1 _5261_/B sky130_fd_sc_hd__or4b_1
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4882_ _5950_/Q _4880_/X _4915_/S vssd1 vssd1 vccd1 vccd1 _4882_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3833_ _3928_/A _5228_/B _3833_/C _3841_/B vssd1 vssd1 vccd1 vccd1 _3834_/B sky130_fd_sc_hd__and4bb_1
X_3764_ _3764_/A vssd1 vssd1 vccd1 vccd1 _5704_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4331__B _4331_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3695_ _3701_/A _3695_/B vssd1 vssd1 vccd1 vccd1 _3696_/A sky130_fd_sc_hd__and2_1
X_5503_ _5529_/A vssd1 vssd1 vccd1 vccd1 _5503_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5434_ _6043_/Q _5439_/B vssd1 vssd1 vccd1 vccd1 _5434_/X sky130_fd_sc_hd__or2_1
XANTENNA__3228__A _6034_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5365_ _5363_/X _5347_/X _5364_/X _5355_/X vssd1 vssd1 vccd1 vccd1 _6021_/D sky130_fd_sc_hd__o211a_1
X_5296_ _5296_/A vssd1 vssd1 vccd1 vccd1 _6009_/D sky130_fd_sc_hd__clkbuf_1
X_4316_ _4316_/A vssd1 vssd1 vccd1 vccd1 _5304_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_59_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4247_ _4249_/B _4228_/X _4246_/Y vssd1 vssd1 vccd1 vccd1 _5805_/D sky130_fd_sc_hd__a21oi_1
XFILLER_87_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4178_ _4178_/A vssd1 vssd1 vccd1 vccd1 _5795_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3129_ _5667_/Q _5713_/Q vssd1 vssd1 vccd1 vccd1 _3129_/X sky130_fd_sc_hd__or2b_1
XFILLER_70_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3410__B _3466_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3908__A2 _4259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5530__A1 _5396_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5353__A input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_43 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3480_ _3480_/A _3480_/B _3480_/C _3486_/A vssd1 vssd1 vccd1 vccd1 _3480_/X sky130_fd_sc_hd__or4_1
XFILLER_6_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2887__A _3839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5521__A1 _5382_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5150_ _5405_/B _5150_/B vssd1 vssd1 vccd1 vccd1 _5168_/B sky130_fd_sc_hd__nor2_1
XFILLER_37_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4101_ _4170_/A vssd1 vssd1 vccd1 vccd1 _4116_/S sky130_fd_sc_hd__buf_2
X_5081_ _5603_/B _5150_/B vssd1 vssd1 vccd1 vccd1 _5100_/B sky130_fd_sc_hd__nor2_1
XFILLER_84_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4032_ _4203_/S vssd1 vssd1 vccd1 vccd1 _4046_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__4607__A _4607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5983_ _5983_/CLK _5983_/D vssd1 vssd1 vccd1 vccd1 _5983_/Q sky130_fd_sc_hd__dfxtp_1
X_4934_ _6038_/Q _4924_/X _4933_/X _4929_/X vssd1 vssd1 vccd1 vccd1 _5912_/D sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_19_wb_clk_i _5836_/CLK vssd1 vssd1 vccd1 vccd1 _6132_/CLK sky130_fd_sc_hd__clkbuf_16
X_4865_ _4819_/X _4863_/X _4864_/X _4824_/X vssd1 vssd1 vccd1 vccd1 _4865_/X sky130_fd_sc_hd__o211a_1
XFILLER_32_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3816_ _3815_/Y _3816_/B vssd1 vssd1 vccd1 vccd1 _5340_/S sky130_fd_sc_hd__and2b_1
X_4796_ _5895_/Q _4756_/X _4794_/X _4795_/X vssd1 vssd1 vccd1 vccd1 _5895_/D sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_13_wb_clk_i_A clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3747_ _3750_/A _3747_/B vssd1 vssd1 vccd1 vccd1 _3748_/A sky130_fd_sc_hd__and2_1
X_3678_ _3582_/A _5681_/Q _3678_/S vssd1 vssd1 vccd1 vccd1 _3679_/B sky130_fd_sc_hd__mux2_1
XANTENNA__5512__A1 _5373_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5417_ _6037_/Q _5417_/B vssd1 vssd1 vccd1 vccd1 _5417_/X sky130_fd_sc_hd__or2_1
X_5348_ _5348_/A vssd1 vssd1 vccd1 vccd1 _5622_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5279_ _5279_/A _5304_/B vssd1 vssd1 vccd1 vccd1 _5280_/A sky130_fd_sc_hd__nand2_1
XFILLER_87_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_52_wb_clk_i_A clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_70_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_proj_example_116 vssd1 vssd1 vccd1 vccd1 user_proj_example_116/HI io_oeb[34]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_105 vssd1 vssd1 vccd1 vccd1 user_proj_example_105/HI io_oeb[23]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_127 vssd1 vssd1 vccd1 vccd1 user_proj_example_127/HI la_data_out[2]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_149 vssd1 vssd1 vccd1 vccd1 user_proj_example_149/HI la_data_out[24]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_138 vssd1 vssd1 vccd1 vccd1 user_proj_example_138/HI la_data_out[13]
+ sky130_fd_sc_hd__conb_1
XFILLER_3_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3331__A _4113_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2980_ _3438_/B _3439_/A _3518_/A vssd1 vssd1 vccd1 vccd1 _3020_/A sky130_fd_sc_hd__a21o_1
XFILLER_61_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5258__A _5258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4650_ _6045_/Q _4584_/X _4610_/X _4649_/X vssd1 vssd1 vccd1 vccd1 _4650_/X sky130_fd_sc_hd__a211o_1
X_3601_ _3601_/A vssd1 vssd1 vccd1 vccd1 _3601_/X sky130_fd_sc_hd__clkbuf_2
Xinput21 la_data_in[47] vssd1 vssd1 vccd1 vccd1 _3582_/A sky130_fd_sc_hd__clkbuf_1
Xinput10 la_data_in[37] vssd1 vssd1 vccd1 vccd1 _5366_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput43 wbs_sel_i[0] vssd1 vssd1 vccd1 vccd1 _3620_/C sky130_fd_sc_hd__clkbuf_1
Xinput32 la_data_in[57] vssd1 vssd1 vccd1 vccd1 _5056_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4581_ _4594_/C vssd1 vssd1 vccd1 vccd1 _4604_/B sky130_fd_sc_hd__clkbuf_2
X_3532_ _5945_/Q _5741_/Q _3561_/B _4568_/B vssd1 vssd1 vccd1 vccd1 _3532_/X sky130_fd_sc_hd__a22o_1
X_3463_ _3481_/B _3463_/B vssd1 vssd1 vccd1 vccd1 _3463_/X sky130_fd_sc_hd__or2_1
X_5202_ _5225_/S vssd1 vssd1 vccd1 vccd1 _5216_/S sky130_fd_sc_hd__clkbuf_2
X_3394_ _3394_/A vssd1 vssd1 vccd1 vccd1 _6131_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5133_ _5056_/X _5125_/X _5132_/X _5130_/X vssd1 vssd1 vccd1 vccd1 _5972_/D sky130_fd_sc_hd__o211a_1
XFILLER_57_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5064_ _5062_/X _5050_/X _5063_/X _5043_/X vssd1 vssd1 vccd1 vccd1 _5950_/D sky130_fd_sc_hd__o211a_1
X_4015_ _2969_/B _3440_/B _4447_/A _4229_/A vssd1 vssd1 vccd1 vccd1 _4016_/B sky130_fd_sc_hd__a211o_1
XFILLER_25_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3241__A _6028_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5966_ _5966_/CLK _5966_/D vssd1 vssd1 vccd1 vccd1 _5966_/Q sky130_fd_sc_hd__dfxtp_1
X_5897_ _6087_/CLK _5897_/D vssd1 vssd1 vccd1 vccd1 _5897_/Q sky130_fd_sc_hd__dfxtp_1
X_4917_ _5970_/Q _4917_/B vssd1 vssd1 vccd1 vccd1 _4917_/X sky130_fd_sc_hd__or2_1
X_4848_ _5997_/Q _5989_/Q _4848_/S vssd1 vssd1 vccd1 vccd1 _4848_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4779_ _4779_/A vssd1 vssd1 vccd1 vccd1 _4821_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_0_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_506 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3151__A _3408_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4472__A1 _5250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4775__A2 _4757_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5078__A _5603_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3735__A0 _5373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3326__A _3326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3061__A _3061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4215__A1 _3880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5820_ _6117_/CLK _5820_/D vssd1 vssd1 vccd1 vccd1 _5820_/Q sky130_fd_sc_hd__dfxtp_1
X_2963_ _5717_/Q _3824_/D vssd1 vssd1 vccd1 vccd1 _3820_/B sky130_fd_sc_hd__nand2_1
X_5751_ _6115_/CLK _5751_/D vssd1 vssd1 vccd1 vccd1 _5751_/Q sky130_fd_sc_hd__dfxtp_1
X_4702_ _6050_/Q _4654_/X _4664_/X _4701_/X vssd1 vssd1 vccd1 vccd1 _4702_/X sky130_fd_sc_hd__a211o_1
X_2894_ _3298_/A vssd1 vssd1 vccd1 vccd1 _3553_/A sky130_fd_sc_hd__clkbuf_2
X_5682_ _5703_/CLK _5682_/D vssd1 vssd1 vccd1 vccd1 _5682_/Q sky130_fd_sc_hd__dfxtp_1
X_4633_ _6043_/Q _4584_/X _4610_/X _4632_/X vssd1 vssd1 vccd1 vccd1 _4633_/X sky130_fd_sc_hd__a211o_1
X_4564_ _5874_/Q _4487_/A _4563_/X _4490_/Y _3723_/C vssd1 vssd1 vccd1 vccd1 _4564_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4620__A _4824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3515_ _4383_/A vssd1 vssd1 vccd1 vccd1 _5278_/A sky130_fd_sc_hd__buf_2
X_4495_ _5860_/Q vssd1 vssd1 vccd1 vccd1 _4518_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3446_ _4470_/C vssd1 vssd1 vccd1 vccd1 _3880_/S sky130_fd_sc_hd__clkbuf_2
X_3377_ _4455_/A _3372_/X _3391_/B _3525_/A vssd1 vssd1 vccd1 vccd1 _3377_/X sky130_fd_sc_hd__o211a_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5116_ _5967_/Q _5116_/B vssd1 vssd1 vccd1 vccd1 _5116_/X sky130_fd_sc_hd__or2_1
X_6096_ _6118_/CLK _6096_/D vssd1 vssd1 vccd1 vccd1 _6096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5047_ _5343_/A _5201_/B vssd1 vssd1 vccd1 vccd1 _5051_/A sky130_fd_sc_hd__nand2_1
XFILLER_72_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_34_wb_clk_i clkbuf_3_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6064_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_53_531 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5949_ _5974_/CLK _5949_/D vssd1 vssd1 vccd1 vccd1 _5949_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3717__B1 _5875_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5626__A _6113_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4390__A0 _6055_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5361__A _6020_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input24_A la_data_in[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4445__A1 _3802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3056__A _3857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3300_ _3300_/A _3300_/B _3300_/C _3299_/X vssd1 vssd1 vccd1 vccd1 _3300_/X sky130_fd_sc_hd__or4b_1
XANTENNA__4920__A2 _5379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4280_ _4280_/A _5813_/Q vssd1 vssd1 vccd1 vccd1 _4281_/D sky130_fd_sc_hd__or2_1
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3231_ _6033_/Q _5934_/Q vssd1 vssd1 vccd1 vccd1 _3231_/Y sky130_fd_sc_hd__nor2_1
X_3162_ _3839_/A _5836_/Q vssd1 vssd1 vccd1 vccd1 _3350_/C sky130_fd_sc_hd__and2_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3093_ _3929_/B vssd1 vssd1 vccd1 vccd1 _3391_/A sky130_fd_sc_hd__buf_2
XFILLER_54_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5803_ _5941_/CLK _5803_/D vssd1 vssd1 vccd1 vccd1 _5803_/Q sky130_fd_sc_hd__dfxtp_1
X_3995_ _3995_/A vssd1 vssd1 vccd1 vccd1 _5735_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2946_ _5327_/A _5309_/A _6010_/Q vssd1 vssd1 vccd1 vccd1 _3400_/B sky130_fd_sc_hd__or3_2
X_5734_ _5808_/CLK _5734_/D vssd1 vssd1 vccd1 vccd1 _5734_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2877_ _3312_/B vssd1 vssd1 vccd1 vccd1 _4464_/B sky130_fd_sc_hd__buf_2
X_5665_ _6112_/CLK _5665_/D vssd1 vssd1 vccd1 vccd1 _5665_/Q sky130_fd_sc_hd__dfxtp_2
X_4616_ _4842_/A vssd1 vssd1 vccd1 vccd1 _5102_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__5446__A _5461_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5596_ _6103_/Q _5599_/B vssd1 vssd1 vccd1 vccd1 _5596_/X sky130_fd_sc_hd__or2_1
X_4547_ _4549_/A _4548_/B _4547_/C vssd1 vssd1 vccd1 vccd1 _5869_/D sky130_fd_sc_hd__nor3_1
XANTENNA__4911__A2 _4706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4478_ _5336_/S _4331_/B _4477_/X _3815_/Y _3274_/B vssd1 vssd1 vccd1 vccd1 _4478_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_1_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3429_ _5323_/B _3429_/B vssd1 vssd1 vccd1 vccd1 _3429_/X sky130_fd_sc_hd__or2_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6079_ _6080_/CLK _6079_/D vssd1 vssd1 vccd1 vccd1 _6079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3780_ _3607_/A _5709_/Q _3780_/S vssd1 vssd1 vccd1 vccd1 _3781_/B sky130_fd_sc_hd__mux2_1
XFILLER_44_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5450_ _5581_/A _5471_/B vssd1 vssd1 vccd1 vccd1 _5467_/B sky130_fd_sc_hd__nor2_1
XANTENNA__4170__A _4170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4401_ _5258_/A _4401_/B vssd1 vssd1 vccd1 vccd1 _5254_/C sky130_fd_sc_hd__and2_1
XFILLER_8_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5381_ _5376_/X _5378_/X _5380_/X _5371_/X vssd1 vssd1 vccd1 vccd1 _6025_/D sky130_fd_sc_hd__o211a_1
X_4332_ _4399_/S vssd1 vssd1 vccd1 vccd1 _4337_/S sky130_fd_sc_hd__dlymetal6s2s_1
X_4263_ _3360_/B _4261_/X _4262_/Y _4231_/A vssd1 vssd1 vccd1 vccd1 _4270_/A sky130_fd_sc_hd__o31a_1
XFILLER_86_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3214_ _3214_/A _3214_/B _3214_/C _3214_/D vssd1 vssd1 vccd1 vccd1 _3215_/C sky130_fd_sc_hd__and4_1
X_6002_ _6002_/CLK _6002_/D vssd1 vssd1 vccd1 vccd1 _6002_/Q sky130_fd_sc_hd__dfxtp_1
X_4194_ _5800_/Q _4193_/X _4200_/S vssd1 vssd1 vccd1 vccd1 _4195_/A sky130_fd_sc_hd__mux2_1
X_3145_ input1/X _3144_/X _5666_/Q vssd1 vssd1 vccd1 vccd1 _3146_/B sky130_fd_sc_hd__mux2_1
XFILLER_27_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3076_ _4240_/B vssd1 vssd1 vccd1 vccd1 _3076_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_49 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3978_ _5730_/Q _3932_/X _3977_/X vssd1 vssd1 vccd1 vccd1 _3979_/B sky130_fd_sc_hd__a21oi_1
X_2929_ _2950_/A _2959_/C _3465_/B _3044_/D vssd1 vssd1 vccd1 vccd1 _3874_/A sky130_fd_sc_hd__or4bb_2
X_5717_ _5796_/CLK _5717_/D vssd1 vssd1 vccd1 vccd1 _5717_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4593__A0 _6089_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5648_ _6135_/Q _5648_/B vssd1 vssd1 vccd1 vccd1 _5648_/X sky130_fd_sc_hd__or2_1
XANTENNA__3408__B _3408_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5542__C1 _5529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5579_ _5579_/A _5601_/B vssd1 vssd1 vccd1 vccd1 _5580_/A sky130_fd_sc_hd__or2_1
XFILLER_77_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3871__A2 _3159_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5086__A _5408_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5300__A2 _5278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output55_A _5882_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput8 la_data_in[35] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_2
XFILLER_76_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2892__B _3494_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4950_ _5918_/Q _4964_/B vssd1 vssd1 vccd1 vccd1 _4953_/B sky130_fd_sc_hd__nand2_1
XANTENNA__4165__A _4182_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3901_ _3901_/A _3901_/B vssd1 vssd1 vccd1 vccd1 _3901_/Y sky130_fd_sc_hd__nand2_1
X_4881_ _4881_/A vssd1 vssd1 vccd1 vccd1 _4915_/S sky130_fd_sc_hd__clkbuf_2
X_3832_ _3832_/A _3903_/A vssd1 vssd1 vccd1 vccd1 _5233_/A sky130_fd_sc_hd__or2_1
XFILLER_20_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3763_ _3768_/A _3763_/B vssd1 vssd1 vccd1 vccd1 _3764_/A sky130_fd_sc_hd__and2_1
X_5502_ _6068_/Q _5505_/B vssd1 vssd1 vccd1 vccd1 _5502_/X sky130_fd_sc_hd__or2_1
XANTENNA__4104__S _4110_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3694_ _3604_/A _5685_/Q _3697_/S vssd1 vssd1 vccd1 vccd1 _3695_/B sky130_fd_sc_hd__mux2_1
X_5433_ _5353_/X _5427_/X _5432_/X _5420_/X vssd1 vssd1 vccd1 vccd1 _6042_/D sky130_fd_sc_hd__o211a_1
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4878__A1 _5981_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5364_ _6021_/Q _5367_/B vssd1 vssd1 vccd1 vccd1 _5364_/X sky130_fd_sc_hd__or2_1
X_4315_ _4315_/A _4315_/B vssd1 vssd1 vccd1 vccd1 _5812_/D sky130_fd_sc_hd__nor2_1
X_5295_ _5295_/A _5295_/B vssd1 vssd1 vccd1 vccd1 _5296_/A sky130_fd_sc_hd__and2_1
X_4246_ _4249_/B _4228_/X _4276_/A vssd1 vssd1 vccd1 vccd1 _4246_/Y sky130_fd_sc_hd__o21bai_1
X_4177_ _5795_/Q _4176_/X _4184_/S vssd1 vssd1 vccd1 vccd1 _4178_/A sky130_fd_sc_hd__mux2_1
X_3128_ _5737_/Q vssd1 vssd1 vccd1 vccd1 _4562_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5055__A1 _5045_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3059_ _3022_/X _3059_/B _3059_/C _3059_/D vssd1 vssd1 vccd1 vccd1 _3059_/X sky130_fd_sc_hd__and4b_1
XFILLER_70_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_42_wb_clk_i_A clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__4802__A1 _6060_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4803__A _5403_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3154__A _4458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4557__A0 _3454_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4100_ _4187_/A vssd1 vssd1 vccd1 vccd1 _4170_/A sky130_fd_sc_hd__clkbuf_2
X_5080_ _5080_/A vssd1 vssd1 vccd1 vccd1 _5080_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3999__A _3999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4031_ _4187_/A vssd1 vssd1 vccd1 vccd1 _4203_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_2_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3835__A2 _3283_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5982_ _5999_/CLK _5982_/D vssd1 vssd1 vccd1 vccd1 _5982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4933_ _5912_/Q _4942_/B vssd1 vssd1 vccd1 vccd1 _4933_/X sky130_fd_sc_hd__or2_1
XFILLER_24_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4623__A _4858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4864_ _5964_/Q _4885_/B vssd1 vssd1 vccd1 vccd1 _4864_/X sky130_fd_sc_hd__or2_1
XFILLER_32_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3815_ _5339_/S _3379_/A _3525_/A vssd1 vssd1 vccd1 vccd1 _3815_/Y sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_59_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6050_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_4795_ _6035_/Q _4744_/X _4745_/X vssd1 vssd1 vccd1 vccd1 _4795_/X sky130_fd_sc_hd__o21a_1
XFILLER_32_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3746_ _5386_/A _5699_/Q _3753_/S vssd1 vssd1 vccd1 vccd1 _3747_/B sky130_fd_sc_hd__mux2_1
XFILLER_9_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3677_ _3677_/A vssd1 vssd1 vccd1 vccd1 _5680_/D sky130_fd_sc_hd__clkbuf_1
X_5416_ _3604_/X _5404_/X _5415_/X _5409_/X vssd1 vssd1 vccd1 vccd1 _6036_/D sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_leaf_9_wb_clk_i_A _5813_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3523__A1 _5278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3523__B2 _3505_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4720__A0 _6100_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5347_ _5354_/B vssd1 vssd1 vccd1 vccd1 _5347_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5278_ _5278_/A _5278_/B _5278_/C _5278_/D vssd1 vssd1 vccd1 vccd1 _5278_/Y sky130_fd_sc_hd__nor4_1
X_4229_ _4229_/A vssd1 vssd1 vccd1 vccd1 _4229_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_231 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_proj_example_117 vssd1 vssd1 vccd1 vccd1 user_proj_example_117/HI io_oeb[35]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_106 vssd1 vssd1 vccd1 vccd1 user_proj_example_106/HI io_oeb[24]
+ sky130_fd_sc_hd__conb_1
XFILLER_11_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xuser_proj_example_128 vssd1 vssd1 vccd1 vccd1 user_proj_example_128/HI la_data_out[3]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_139 vssd1 vssd1 vccd1 vccd1 user_proj_example_139/HI la_data_out[14]
+ sky130_fd_sc_hd__conb_1
XANTENNA__2988__A _3518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5364__A _6021_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3514__A1 _3135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5258__B _5258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4580_ _4580_/A _3564_/B vssd1 vssd1 vccd1 vccd1 _4594_/C sky130_fd_sc_hd__or2b_1
Xinput22 la_data_in[48] vssd1 vssd1 vccd1 vccd1 _3587_/A sky130_fd_sc_hd__clkbuf_1
Xinput11 la_data_in[38] vssd1 vssd1 vccd1 vccd1 _5369_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3600_ _3598_/X _3592_/X _3599_/X _3585_/X vssd1 vssd1 vccd1 vccd1 _5659_/D sky130_fd_sc_hd__o211a_1
X_3531_ _5739_/Q vssd1 vssd1 vccd1 vccd1 _4568_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xinput44 wbs_sel_i[1] vssd1 vssd1 vccd1 vccd1 _3572_/C sky130_fd_sc_hd__clkbuf_1
Xinput33 la_data_in[58] vssd1 vssd1 vccd1 vccd1 _5059_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2898__A _3553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3462_ _3466_/A _3480_/C _3462_/C vssd1 vssd1 vccd1 vccd1 _3462_/X sky130_fd_sc_hd__or3_1
X_3393_ _3632_/A _3393_/B vssd1 vssd1 vccd1 vccd1 _3394_/A sky130_fd_sc_hd__and2_1
X_5201_ _5201_/A _5201_/B vssd1 vssd1 vccd1 vccd1 _5225_/S sky130_fd_sc_hd__nand2_2
XFILLER_69_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5132_ _5972_/Q _5138_/B vssd1 vssd1 vccd1 vccd1 _5132_/X sky130_fd_sc_hd__or2_1
XFILLER_84_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5063_ _5950_/Q _5066_/B vssd1 vssd1 vccd1 vccd1 _5063_/X sky130_fd_sc_hd__or2_1
XANTENNA__4618__A _6066_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4014_ _5247_/A vssd1 vssd1 vccd1 vccd1 _4014_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5965_ _5983_/CLK _5965_/D vssd1 vssd1 vccd1 vccd1 _5965_/Q sky130_fd_sc_hd__dfxtp_1
X_5896_ _6088_/CLK _5896_/D vssd1 vssd1 vccd1 vccd1 _5896_/Q sky130_fd_sc_hd__dfxtp_1
X_4916_ _5962_/Q _4915_/X _4916_/S vssd1 vssd1 vccd1 vccd1 _4916_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4847_ _5900_/Q _4807_/X _4845_/X _4846_/X vssd1 vssd1 vccd1 vccd1 _5900_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4778_ _5706_/Q _5683_/Q _4797_/S vssd1 vssd1 vccd1 vccd1 _4778_/X sky130_fd_sc_hd__mux2_1
X_3729_ _3732_/A _3729_/B vssd1 vssd1 vccd1 vccd1 _3730_/A sky130_fd_sc_hd__and2_1
XANTENNA__5497__A1 _5342_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_518 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5421__A1 _3611_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5185__A0 _5062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_4_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6118_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4202__S _4554_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4215__A2 _3432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2962_ _2994_/B vssd1 vssd1 vccd1 vccd1 _3824_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_5750_ _5796_/CLK _5750_/D vssd1 vssd1 vccd1 vccd1 _5750_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5681_ _5703_/CLK _5681_/D vssd1 vssd1 vccd1 vccd1 _5681_/Q sky130_fd_sc_hd__dfxtp_1
X_4701_ _4665_/X _4699_/X _4700_/X _4670_/X vssd1 vssd1 vccd1 vccd1 _4701_/X sky130_fd_sc_hd__o211a_1
X_2893_ hold1/A vssd1 vssd1 vccd1 vccd1 _3298_/A sky130_fd_sc_hd__inv_2
XANTENNA__5176__A0 _5045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4632_ _4611_/X _4630_/X _4631_/X _4620_/X vssd1 vssd1 vccd1 vccd1 _4632_/X sky130_fd_sc_hd__o211a_1
XFILLER_30_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4563_ _4562_/A _5737_/Q _3553_/X vssd1 vssd1 vccd1 vccd1 _4563_/X sky130_fd_sc_hd__o21ba_1
X_4494_ _4489_/Y _4493_/X _3999_/A vssd1 vssd1 vccd1 vccd1 _5859_/D sky130_fd_sc_hd__a21oi_1
X_3514_ _3135_/A _3350_/A _5269_/B vssd1 vssd1 vccd1 vccd1 _3514_/X sky130_fd_sc_hd__a21o_1
XFILLER_89_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3445_ _2955_/C _3443_/X _3444_/X _3047_/X vssd1 vssd1 vccd1 vccd1 _3452_/A sky130_fd_sc_hd__a22o_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3376_ _3410_/C vssd1 vssd1 vccd1 vccd1 _3525_/A sky130_fd_sc_hd__buf_2
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5115_ _5062_/X _5104_/X _5113_/X _5114_/X vssd1 vssd1 vccd1 vccd1 _5966_/D sky130_fd_sc_hd__o211a_1
X_6095_ _6118_/CLK _6095_/D vssd1 vssd1 vccd1 vccd1 _6095_/Q sky130_fd_sc_hd__dfxtp_1
X_5046_ _5046_/A _5046_/B _5046_/C vssd1 vssd1 vccd1 vccd1 _5201_/B sky130_fd_sc_hd__and3_2
XFILLER_84_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5651__A1 _5389_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4083__A _4203_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5948_ _5974_/CLK _5948_/D vssd1 vssd1 vccd1 vccd1 _5948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5879_ _6024_/CLK _5879_/D vssd1 vssd1 vccd1 vccd1 _5879_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3717__A1 _4575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5642__A _6120_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2985__B _4218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input17_A la_data_in[43] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3230_ _6033_/Q _5934_/Q vssd1 vssd1 vccd1 vccd1 _3230_/X sky130_fd_sc_hd__and2_1
X_3161_ _3161_/A vssd1 vssd1 vccd1 vccd1 _3161_/X sky130_fd_sc_hd__clkbuf_2
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3072__A _3824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3892__B1 _5768_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3092_ _3423_/A _3423_/B _3092_/C _3272_/B vssd1 vssd1 vccd1 vccd1 _3092_/X sky130_fd_sc_hd__or4_1
XFILLER_66_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3644__A0 _5366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4107__S _4110_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5802_ _5929_/CLK _5802_/D vssd1 vssd1 vccd1 vccd1 _5802_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3994_ _3994_/A _3994_/B vssd1 vssd1 vccd1 vccd1 _3995_/A sky130_fd_sc_hd__and2_1
XFILLER_22_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5733_ _5808_/CLK _5733_/D vssd1 vssd1 vccd1 vccd1 _5733_/Q sky130_fd_sc_hd__dfxtp_1
X_2945_ _4218_/B vssd1 vssd1 vccd1 vccd1 _5247_/B sky130_fd_sc_hd__clkbuf_2
X_2876_ _2950_/B vssd1 vssd1 vccd1 vccd1 _2944_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__4631__A _6067_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5664_ _6112_/CLK _5664_/D vssd1 vssd1 vccd1 vccd1 _5664_/Q sky130_fd_sc_hd__dfxtp_1
X_5595_ _5396_/X _5580_/A _5594_/X _5586_/X vssd1 vssd1 vccd1 vccd1 _6102_/D sky130_fd_sc_hd__o211a_1
X_4615_ _6090_/Q _4613_/X _5603_/B vssd1 vssd1 vccd1 vccd1 _4615_/X sky130_fd_sc_hd__mux2_1
X_4546_ _4545_/B _4545_/C _4545_/A vssd1 vssd1 vccd1 vccd1 _4547_/C sky130_fd_sc_hd__a21oi_1
X_4477_ _3161_/X _3274_/B _3260_/X _5716_/Q vssd1 vssd1 vccd1 vccd1 _4477_/X sky130_fd_sc_hd__a31o_1
XFILLER_89_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3428_ _3428_/A _3428_/B _2863_/X vssd1 vssd1 vccd1 vccd1 _3428_/X sky130_fd_sc_hd__or3b_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3359_ _5247_/A _5717_/Q vssd1 vssd1 vccd1 vccd1 _3821_/C sky130_fd_sc_hd__nor2_2
XANTENNA__4078__A _4095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input9_A la_data_in[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6078_ _6080_/CLK _6078_/D vssd1 vssd1 vccd1 vccd1 _6078_/Q sky130_fd_sc_hd__dfxtp_1
X_5029_ _5029_/A _5029_/B vssd1 vssd1 vccd1 vccd1 _5940_/D sky130_fd_sc_hd__nor2_1
XANTENNA__3635__A0 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5637__A _6118_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_443 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4716__A _4716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4400_ _4400_/A vssd1 vssd1 vccd1 vccd1 _5836_/D sky130_fd_sc_hd__clkbuf_1
X_5380_ _6025_/Q _5399_/B vssd1 vssd1 vccd1 vccd1 _5380_/X sky130_fd_sc_hd__or2_1
X_4331_ _4450_/B _4331_/B vssd1 vssd1 vccd1 vccd1 _4399_/S sky130_fd_sc_hd__nand2_2
XFILLER_5_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4262_ _3435_/A _2975_/Y _2982_/B vssd1 vssd1 vccd1 vccd1 _4262_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_4_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3213_ _6023_/Q _3198_/Y _5012_/A _6017_/Q _3212_/X vssd1 vssd1 vccd1 vccd1 _3214_/D
+ sky130_fd_sc_hd__a221oi_1
X_6001_ _6002_/CLK _6001_/D vssd1 vssd1 vccd1 vccd1 _6001_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4193_ _5950_/Q _5799_/Q _4196_/S vssd1 vssd1 vccd1 vccd1 _4193_/X sky130_fd_sc_hd__mux2_1
X_3144_ _5874_/Q _5849_/Q vssd1 vssd1 vccd1 vccd1 _3144_/X sky130_fd_sc_hd__xor2_1
XFILLER_67_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3075_ _3349_/C _3075_/B vssd1 vssd1 vccd1 vccd1 _4240_/B sky130_fd_sc_hd__or2_1
XFILLER_82_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_32_wb_clk_i_A _5836_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3977_ _5729_/Q _3941_/X _3953_/X _3976_/Y vssd1 vssd1 vccd1 vccd1 _3977_/X sky130_fd_sc_hd__o211a_1
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2928_ _3448_/A _2928_/B vssd1 vssd1 vccd1 vccd1 _2928_/Y sky130_fd_sc_hd__nor2_1
X_5716_ _6018_/CLK _5716_/D vssd1 vssd1 vccd1 vccd1 _5716_/Q sky130_fd_sc_hd__dfxtp_1
X_2859_ _6006_/Q vssd1 vssd1 vccd1 vccd1 _5277_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_5647_ _5382_/X _3576_/X _5646_/X _5638_/X vssd1 vssd1 vccd1 vccd1 _6134_/D sky130_fd_sc_hd__o211a_1
X_5578_ _5373_/X _5559_/A _5577_/X _5571_/X vssd1 vssd1 vccd1 vccd1 _6096_/D sky130_fd_sc_hd__o211a_1
X_4529_ _4529_/A _4529_/B vssd1 vssd1 vccd1 vccd1 _4538_/B sky130_fd_sc_hd__and2_1
XANTENNA__3705__A _3732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5058__C1 _5043_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4536__A _4970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5367__A _6022_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4336__B2 _6067_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput9 la_data_in[36] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_91_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3900_ _3821_/A _3821_/C _3899_/Y _3886_/Y vssd1 vssd1 vccd1 vccd1 _3902_/C sky130_fd_sc_hd__a31o_1
XFILLER_51_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4880_ _6000_/Q _5992_/Q _4898_/S vssd1 vssd1 vccd1 vccd1 _4880_/X sky130_fd_sc_hd__mux2_1
X_3831_ _5250_/A _6121_/Q vssd1 vssd1 vccd1 vccd1 _3903_/A sky130_fd_sc_hd__nor2_1
X_3762_ _3582_/A _5704_/Q _3762_/S vssd1 vssd1 vccd1 vccd1 _3763_/B sky130_fd_sc_hd__mux2_1
X_5501_ _5357_/X _5493_/X _5500_/X _5488_/X vssd1 vssd1 vccd1 vccd1 _6067_/D sky130_fd_sc_hd__o211a_1
X_3693_ _3693_/A vssd1 vssd1 vccd1 vccd1 _5684_/D sky130_fd_sc_hd__clkbuf_1
X_5432_ _6042_/Q _5439_/B vssd1 vssd1 vccd1 vccd1 _5432_/X sky130_fd_sc_hd__or2_1
X_5363_ input9/X vssd1 vssd1 vccd1 vccd1 _5363_/X sky130_fd_sc_hd__clkbuf_2
X_4314_ _5812_/Q _4314_/B vssd1 vssd1 vccd1 vccd1 _4315_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__3525__A _3525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5294_ _5297_/B _5293_/X _5294_/S vssd1 vssd1 vccd1 vccd1 _5295_/B sky130_fd_sc_hd__mux2_1
X_4245_ _4233_/X _4228_/X _4244_/Y _3408_/B vssd1 vssd1 vccd1 vccd1 _4276_/A sky130_fd_sc_hd__a31o_1
X_4176_ _5663_/Q _5794_/Q _4179_/S vssd1 vssd1 vccd1 vccd1 _4176_/X sky130_fd_sc_hd__mux2_1
X_3127_ _3127_/A _3127_/B _3127_/C vssd1 vssd1 vccd1 vccd1 _6128_/D sky130_fd_sc_hd__nand3_1
XFILLER_55_413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4246__B1_N _4276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3260__A _4322_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3058_ _3058_/A _3058_/B vssd1 vssd1 vccd1 vccd1 _3059_/D sky130_fd_sc_hd__or2_1
XFILLER_82_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4802__A2 _4757_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4318__A1 _5301_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3170__A _3632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3057__A1 _3375_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3345__A _3841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4030_ _6094_/Q _2858_/A _5752_/Q _4017_/X vssd1 vssd1 vccd1 vccd1 _4030_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5560__A _5603_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4245__B1 _3408_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5981_ _5983_/CLK _5981_/D vssd1 vssd1 vccd1 vccd1 _5981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4932_ _6037_/Q _4924_/X _4931_/Y _4929_/X vssd1 vssd1 vccd1 vccd1 _5911_/D sky130_fd_sc_hd__o211a_1
XANTENNA__4796__A1 _5895_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4260__A3 _3440_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4863_ _5956_/Q _4862_/X _4873_/S vssd1 vssd1 vccd1 vccd1 _4863_/X sky130_fd_sc_hd__mux2_1
X_3814_ _4237_/C _3814_/B _3814_/C vssd1 vssd1 vccd1 vccd1 _3816_/B sky130_fd_sc_hd__or3_1
X_4794_ _6059_/Q _4757_/X _4767_/X _4793_/X vssd1 vssd1 vccd1 vccd1 _4794_/X sky130_fd_sc_hd__a211o_1
X_3745_ _3745_/A vssd1 vssd1 vccd1 vccd1 _5698_/D sky130_fd_sc_hd__clkbuf_1
X_3676_ _3684_/A _3676_/B vssd1 vssd1 vccd1 vccd1 _3677_/A sky130_fd_sc_hd__and2_1
X_5415_ _6036_/Q _5417_/B vssd1 vssd1 vccd1 vccd1 _5415_/X sky130_fd_sc_hd__or2_1
XANTENNA__3255__A _3668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_28_wb_clk_i clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5914_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_5346_ _5346_/A vssd1 vssd1 vccd1 vccd1 _5354_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5277_ _5277_/A _5277_/B _5277_/C vssd1 vssd1 vccd1 vccd1 _5297_/C sky130_fd_sc_hd__and3_1
X_4228_ _4249_/C vssd1 vssd1 vccd1 vccd1 _4228_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_75_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4159_ _5658_/Q _3480_/B _4162_/S vssd1 vssd1 vccd1 vccd1 _4159_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5433__C1 _5420_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xuser_proj_example_118 vssd1 vssd1 vccd1 vccd1 user_proj_example_118/HI io_oeb[36]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_107 vssd1 vssd1 vccd1 vccd1 user_proj_example_107/HI io_oeb[25]
+ sky130_fd_sc_hd__conb_1
XANTENNA__3211__B2 _6017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xuser_proj_example_129 vssd1 vssd1 vccd1 vccd1 user_proj_example_129/HI la_data_out[4]
+ sky130_fd_sc_hd__conb_1
XFILLER_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input47_A wbs_stb_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5380__A _6025_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput12 la_data_in[39] vssd1 vssd1 vccd1 vccd1 _5373_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3530_ _5857_/Q _3529_/Y _4480_/A vssd1 vssd1 vccd1 vccd1 _3561_/B sky130_fd_sc_hd__o21ai_1
Xinput23 la_data_in[49] vssd1 vssd1 vccd1 vccd1 _3598_/A sky130_fd_sc_hd__clkbuf_1
Xinput45 wbs_sel_i[2] vssd1 vssd1 vccd1 vccd1 _3588_/B sky130_fd_sc_hd__clkbuf_1
Xinput34 la_data_in[59] vssd1 vssd1 vccd1 vccd1 _5062_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2898__B _3469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3461_ _3854_/A vssd1 vssd1 vccd1 vccd1 _3480_/C sky130_fd_sc_hd__clkbuf_2
X_3392_ _5249_/A _3522_/A _3390_/Y _3391_/Y _4455_/A vssd1 vssd1 vccd1 vccd1 _3393_/B
+ sky130_fd_sc_hd__a32o_1
X_5200_ _5200_/A vssd1 vssd1 vccd1 vccd1 _5996_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5131_ _5045_/X _5125_/X _5129_/X _5130_/X vssd1 vssd1 vccd1 vccd1 _5971_/D sky130_fd_sc_hd__o211a_1
X_5062_ _5062_/A vssd1 vssd1 vccd1 vccd1 _5062_/X sky130_fd_sc_hd__clkbuf_2
X_4013_ _6089_/Q _3061_/A _4028_/S _4012_/X vssd1 vssd1 vccd1 vccd1 _5748_/D sky130_fd_sc_hd__a31o_1
XANTENNA__4618__B _5537_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5964_ _5983_/CLK _5964_/D vssd1 vssd1 vccd1 vccd1 _5964_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3441__A1 _3326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5895_ _6088_/CLK _5895_/D vssd1 vssd1 vccd1 vccd1 _5895_/Q sky130_fd_sc_hd__dfxtp_1
X_4915_ _5954_/Q _4914_/X _4915_/S vssd1 vssd1 vccd1 vccd1 _4915_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4846_ _6040_/Q _4803_/X _4804_/X vssd1 vssd1 vccd1 vccd1 _4846_/X sky130_fd_sc_hd__o21a_1
XANTENNA__4941__A1 _5979_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5465__A _6055_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4777_ _5893_/Q _4756_/X _4775_/X _4776_/X vssd1 vssd1 vccd1 vccd1 _5893_/D sky130_fd_sc_hd__a22o_1
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3728_ _5366_/A _5694_/Q _3735_/S vssd1 vssd1 vccd1 vccd1 _3729_/B sky130_fd_sc_hd__mux2_1
X_3659_ _5382_/A _5675_/Q _3669_/S vssd1 vssd1 vccd1 vccd1 _3660_/B sky130_fd_sc_hd__mux2_1
X_5329_ _5262_/X _5326_/X _5328_/X _3547_/A vssd1 vssd1 vccd1 vccd1 _5329_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3833__A_N _3928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3713__A _3794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3432__B _3432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4932__A1 _6037_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4438__B _4438_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2961_ _5812_/Q _5811_/Q _5810_/Q _5809_/Q vssd1 vssd1 vccd1 vccd1 _2994_/B sky130_fd_sc_hd__and4bb_1
X_5680_ _5703_/CLK _5680_/D vssd1 vssd1 vccd1 vccd1 _5680_/Q sky130_fd_sc_hd__dfxtp_1
X_4700_ _6074_/Q _4732_/B vssd1 vssd1 vccd1 vccd1 _4700_/X sky130_fd_sc_hd__or2_1
X_2892_ _3480_/B _3494_/B _3304_/B vssd1 vssd1 vccd1 vccd1 _2892_/X sky130_fd_sc_hd__and3_1
XFILLER_30_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4631_ _6067_/Q _5537_/B vssd1 vssd1 vccd1 vccd1 _4631_/X sky130_fd_sc_hd__or2_1
XANTENNA__4901__B _4917_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4562_ _4562_/A _4562_/B _5847_/Q vssd1 vssd1 vccd1 vccd1 _4562_/X sky130_fd_sc_hd__or3_1
X_4493_ _4562_/B _4490_/Y _4489_/B _3538_/Y vssd1 vssd1 vccd1 vccd1 _4493_/X sky130_fd_sc_hd__a211o_1
X_3513_ _4383_/A _3513_/B vssd1 vssd1 vccd1 vccd1 _5269_/B sky130_fd_sc_hd__and2_1
X_3444_ _3858_/A _3035_/C _3042_/X _3440_/B _3046_/Y vssd1 vssd1 vccd1 vccd1 _3444_/X
+ sky130_fd_sc_hd__a41o_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3375_ _3553_/A _3375_/B vssd1 vssd1 vccd1 vccd1 _3410_/C sky130_fd_sc_hd__nor2_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5114_ _5141_/A vssd1 vssd1 vccd1 vccd1 _5114_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6094_ _6118_/CLK _6094_/D vssd1 vssd1 vccd1 vccd1 _6094_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5045_ _5045_/A vssd1 vssd1 vccd1 vccd1 _5045_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_72_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5947_ _6040_/CLK _5947_/D vssd1 vssd1 vccd1 vccd1 _5947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5878_ _6108_/CLK _5878_/D vssd1 vssd1 vccd1 vccd1 _5878_/Q sky130_fd_sc_hd__dfxtp_1
X_4829_ _5711_/Q _5688_/Q _4848_/S vssd1 vssd1 vccd1 vccd1 _4829_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_43_wb_clk_i clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6002_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__3708__A _3732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4539__A _4970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3618__A _5665_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3160_ _5241_/B _3257_/A vssd1 vssd1 vccd1 vccd1 _3484_/B sky130_fd_sc_hd__nand2_4
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__dlygate4sd3_1
X_3091_ _3411_/B vssd1 vssd1 vccd1 vccd1 _3423_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_clkbuf_leaf_22_wb_clk_i_A clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_81_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4841__A0 _6112_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5801_ _5929_/CLK _5801_/D vssd1 vssd1 vccd1 vccd1 _5801_/Q sky130_fd_sc_hd__dfxtp_1
X_5732_ _5808_/CLK _5732_/D vssd1 vssd1 vccd1 vccd1 _5732_/Q sky130_fd_sc_hd__dfxtp_1
X_3993_ _5735_/Q _3964_/A _3953_/A _5734_/Q vssd1 vssd1 vccd1 vccd1 _3994_/B sky130_fd_sc_hd__a22o_1
XFILLER_62_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2944_ _3321_/A _2944_/B _4464_/B _3465_/C vssd1 vssd1 vccd1 vccd1 _4218_/B sky130_fd_sc_hd__nor4b_4
X_2875_ _4281_/C vssd1 vssd1 vccd1 vccd1 _3853_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4631__B _5537_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5663_ _6109_/CLK _5663_/D vssd1 vssd1 vccd1 vccd1 _5663_/Q sky130_fd_sc_hd__dfxtp_1
X_5594_ _6102_/Q _5599_/B vssd1 vssd1 vccd1 vccd1 _5594_/X sky130_fd_sc_hd__or2_1
X_4614_ _4883_/A vssd1 vssd1 vccd1 vccd1 _5603_/B sky130_fd_sc_hd__buf_2
X_4545_ _4545_/A _4545_/B _4545_/C vssd1 vssd1 vccd1 vccd1 _4548_/B sky130_fd_sc_hd__and3_1
X_4476_ _4476_/A vssd1 vssd1 vccd1 vccd1 _5851_/D sky130_fd_sc_hd__clkbuf_1
X_3427_ _3460_/A _5320_/A _3427_/C vssd1 vssd1 vccd1 vccd1 _3427_/X sky130_fd_sc_hd__or3_1
XANTENNA_clkbuf_leaf_61_wb_clk_i_A clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__3332__B1 _3331_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3358_ _3357_/X _3898_/A _3341_/B _3256_/A _3350_/A vssd1 vssd1 vccd1 vccd1 _3520_/B
+ sky130_fd_sc_hd__o2111a_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3289_ _3849_/A vssd1 vssd1 vccd1 vccd1 _3897_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6077_ _6077_/CLK _6077_/D vssd1 vssd1 vccd1 vccd1 _6077_/Q sky130_fd_sc_hd__dfxtp_1
X_5028_ _5940_/Q _5030_/C _5020_/X vssd1 vssd1 vccd1 vccd1 _5029_/B sky130_fd_sc_hd__o21ai_1
XFILLER_57_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5388__A1 _5386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_455 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3551__A_N _5667_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_499 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4330_ _4288_/Y _4328_/X _4329_/Y _2955_/C vssd1 vssd1 vccd1 vccd1 _5813_/D sky130_fd_sc_hd__o2bb2a_1
XFILLER_4_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4261_ _3880_/S _4258_/X _4259_/Y _4260_/X vssd1 vssd1 vccd1 vccd1 _4261_/X sky130_fd_sc_hd__o31a_1
XFILLER_5_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3212_ _6021_/Q _5940_/Q vssd1 vssd1 vccd1 vccd1 _3212_/X sky130_fd_sc_hd__xor2_1
X_6000_ _6002_/CLK _6000_/D vssd1 vssd1 vccd1 vccd1 _6000_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4192_ _4192_/A vssd1 vssd1 vccd1 vccd1 _5799_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3143_ _5849_/Q vssd1 vssd1 vccd1 vccd1 _4567_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_82_425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3074_ _3873_/A _3092_/C vssd1 vssd1 vccd1 vccd1 _3075_/B sky130_fd_sc_hd__nor2_1
XFILLER_67_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4290__A1 _3802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3976_ _5729_/Q _3983_/B vssd1 vssd1 vccd1 vccd1 _3976_/Y sky130_fd_sc_hd__nand2_1
X_2927_ _4255_/A _2863_/A _3058_/A _3015_/A vssd1 vssd1 vccd1 vccd1 _2928_/B sky130_fd_sc_hd__o211a_1
X_5715_ _6018_/CLK _5715_/D vssd1 vssd1 vccd1 vccd1 _5715_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5646_ _6134_/Q _5648_/B vssd1 vssd1 vccd1 vccd1 _5646_/X sky130_fd_sc_hd__or2_1
X_2858_ _2858_/A vssd1 vssd1 vccd1 vccd1 _3061_/A sky130_fd_sc_hd__clkbuf_2
X_5577_ _6096_/Q _5577_/B vssd1 vssd1 vccd1 vccd1 _5577_/X sky130_fd_sc_hd__or2_1
X_4528_ _4567_/A _3544_/B _3556_/B vssd1 vssd1 vccd1 vccd1 _4529_/B sky130_fd_sc_hd__o21a_1
XFILLER_2_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4459_ _5408_/A vssd1 vssd1 vccd1 vccd1 _5067_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6129_ _6130_/CLK _6129_/D vssd1 vssd1 vccd1 vccd1 _6129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_355 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5558__A _5601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3830_ _4471_/A _3830_/B vssd1 vssd1 vccd1 vccd1 _3832_/A sky130_fd_sc_hd__nor2_1
XFILLER_32_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3761_ _3761_/A vssd1 vssd1 vccd1 vccd1 _5703_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3078__A _5255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5500_ _6067_/Q _5505_/B vssd1 vssd1 vccd1 vccd1 _5500_/X sky130_fd_sc_hd__or2_1
XANTENNA__3509__C _3954_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4980__C1 _3255_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3692_ _3701_/A _3692_/B vssd1 vssd1 vccd1 vccd1 _3693_/A sky130_fd_sc_hd__and2_1
X_5431_ _5342_/X _5427_/X _5430_/X _5420_/X vssd1 vssd1 vccd1 vccd1 _6041_/D sky130_fd_sc_hd__o211a_1
X_5362_ _5360_/X _5347_/X _5361_/X _5355_/X vssd1 vssd1 vccd1 vccd1 _6020_/D sky130_fd_sc_hd__o211a_1
X_4313_ _5811_/Q _5810_/Q _4313_/C vssd1 vssd1 vccd1 vccd1 _4314_/B sky130_fd_sc_hd__and3_1
X_5293_ _5323_/A _5288_/D _5287_/X _5292_/X vssd1 vssd1 vccd1 vccd1 _5293_/X sky130_fd_sc_hd__a31o_1
XFILLER_87_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4244_ _4244_/A vssd1 vssd1 vccd1 vccd1 _4244_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4175_ _4175_/A vssd1 vssd1 vccd1 vccd1 _5794_/D sky130_fd_sc_hd__clkbuf_1
X_3126_ _3423_/C _3086_/X _3092_/X _3123_/Y _3547_/A vssd1 vssd1 vccd1 vccd1 _3127_/C
+ sky130_fd_sc_hd__o32a_1
XFILLER_55_425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3057_ _3375_/B _3427_/C _3841_/C _3055_/X _3460_/C vssd1 vssd1 vccd1 vccd1 _3058_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_50_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3959_ _3979_/A _3959_/B vssd1 vssd1 vccd1 vccd1 _5725_/D sky130_fd_sc_hd__nor2_1
X_5629_ _6114_/Q _5635_/B vssd1 vssd1 vccd1 vccd1 _5629_/X sky130_fd_sc_hd__or2_1
XFILLER_2_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5203__A0 _5045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5506__A1 _5363_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3517__B1 _3071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3626__A _5343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output60_A _5887_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5980_ _5983_/CLK _5980_/D vssd1 vssd1 vccd1 vccd1 _5980_/Q sky130_fd_sc_hd__dfxtp_1
X_4931_ _4931_/A _4944_/B vssd1 vssd1 vccd1 vccd1 _4931_/Y sky130_fd_sc_hd__nand2_1
XFILLER_52_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4862_ _5948_/Q _4861_/X _4872_/S vssd1 vssd1 vccd1 vccd1 _4862_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3813_ _3813_/A vssd1 vssd1 vccd1 vccd1 _5715_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4793_ _4768_/X _4790_/X _4792_/X _4773_/X vssd1 vssd1 vccd1 vccd1 _4793_/X sky130_fd_sc_hd__o211a_1
X_3744_ _3750_/A _3744_/B vssd1 vssd1 vccd1 vccd1 _3745_/A sky130_fd_sc_hd__and2_1
XFILLER_20_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3675_ _3563_/A _5680_/Q _3678_/S vssd1 vssd1 vccd1 vccd1 _3676_/B sky130_fd_sc_hd__mux2_1
X_5414_ _3601_/X _5404_/X _5413_/X _5409_/X vssd1 vssd1 vccd1 vccd1 _6035_/D sky130_fd_sc_hd__o211a_1
XFILLER_87_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5345_ _5345_/A _5624_/B vssd1 vssd1 vccd1 vccd1 _5346_/A sky130_fd_sc_hd__or2_1
X_5276_ _5277_/B _5243_/A _5262_/X _5281_/A vssd1 vssd1 vccd1 vccd1 _5284_/B sky130_fd_sc_hd__a31oi_1
XFILLER_87_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4227_ _4213_/X _4227_/B _4227_/C vssd1 vssd1 vccd1 vccd1 _4249_/C sky130_fd_sc_hd__and3b_1
XFILLER_28_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4158_ _4158_/A vssd1 vssd1 vccd1 vccd1 _5789_/D sky130_fd_sc_hd__clkbuf_1
X_3109_ _5234_/A vssd1 vssd1 vccd1 vccd1 _3820_/A sky130_fd_sc_hd__clkbuf_2
X_4089_ _5956_/Q _5769_/Q _4092_/S vssd1 vssd1 vccd1 vccd1 _4089_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_proj_example_108 vssd1 vssd1 vccd1 vccd1 user_proj_example_108/HI io_oeb[26]
+ sky130_fd_sc_hd__conb_1
XFILLER_11_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_proj_example_119 vssd1 vssd1 vccd1 vccd1 user_proj_example_119/HI io_oeb[37]
+ sky130_fd_sc_hd__conb_1
XANTENNA__4041__S _4041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3880__S _3880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4277__A _5736_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_439 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput13 la_data_in[3] vssd1 vssd1 vccd1 vccd1 _3711_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput46 wbs_sel_i[3] vssd1 vssd1 vccd1 vccd1 _5046_/C sky130_fd_sc_hd__clkbuf_1
Xinput35 la_data_in[5] vssd1 vssd1 vccd1 vccd1 _5046_/A sky130_fd_sc_hd__clkbuf_1
Xinput24 la_data_in[4] vssd1 vssd1 vccd1 vccd1 _4580_/A sky130_fd_sc_hd__clkbuf_1
X_3460_ _3460_/A _5320_/A _3460_/C _3460_/D vssd1 vssd1 vccd1 vccd1 _3460_/X sky130_fd_sc_hd__or4_1
X_3391_ _3391_/A _3391_/B vssd1 vssd1 vccd1 vccd1 _3391_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5571__A _5597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5130_ _5141_/A vssd1 vssd1 vccd1 vccd1 _5130_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5061_ _5059_/X _5050_/X _5060_/X _5043_/X vssd1 vssd1 vccd1 vccd1 _5949_/D sky130_fd_sc_hd__o211a_1
XFILLER_84_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3091__A _3411_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4012_ _4010_/A _4473_/B _5748_/Q vssd1 vssd1 vccd1 vccd1 _4012_/X sky130_fd_sc_hd__o21a_1
XFILLER_77_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5963_ _5975_/CLK _5963_/D vssd1 vssd1 vccd1 vccd1 _5963_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4914_ _6004_/Q _5996_/Q _4914_/S vssd1 vssd1 vccd1 vccd1 _4914_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5894_ _6085_/CLK _5894_/D vssd1 vssd1 vccd1 vccd1 _5894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4845_ _6064_/Q _4808_/X _4818_/X _4844_/X vssd1 vssd1 vccd1 vccd1 _4845_/X sky130_fd_sc_hd__a211o_1
XFILLER_32_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4926__C1 _4460_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4776_ _6033_/Q _4744_/X _4745_/X vssd1 vssd1 vccd1 vccd1 _4776_/X sky130_fd_sc_hd__o21a_1
X_3727_ _3727_/A vssd1 vssd1 vccd1 vccd1 _5693_/D sky130_fd_sc_hd__clkbuf_1
X_3658_ _3658_/A vssd1 vssd1 vccd1 vccd1 _5674_/D sky130_fd_sc_hd__clkbuf_1
X_3589_ _5343_/A _3765_/A vssd1 vssd1 vccd1 vccd1 _3593_/A sky130_fd_sc_hd__nand2_1
X_5328_ _3491_/X _5257_/Y _5327_/X _5322_/X _5323_/X vssd1 vssd1 vccd1 vccd1 _5328_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_87_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5481__A _6060_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5259_ _5255_/X _5257_/Y _5258_/Y _5243_/B vssd1 vssd1 vccd1 vccd1 _5259_/X sky130_fd_sc_hd__a31o_1
XFILLER_28_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3499__A2 _3505_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5391__A _5391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4696__A1 _5885_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_12_wb_clk_i_A _5813_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_328 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2960_ _3518_/A _3283_/B vssd1 vssd1 vccd1 vccd1 _3440_/A sky130_fd_sc_hd__nor2_1
X_2891_ _3837_/A vssd1 vssd1 vccd1 vccd1 _3494_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_30_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4630_ _6091_/Q _4628_/X _4668_/S vssd1 vssd1 vccd1 vccd1 _4630_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4561_ _5873_/Q _3551_/X _3245_/X vssd1 vssd1 vccd1 vccd1 _5873_/D sky130_fd_sc_hd__o21a_1
X_4492_ _4489_/Y _4491_/X _5171_/A vssd1 vssd1 vccd1 vccd1 _5858_/D sky130_fd_sc_hd__a21o_1
X_3512_ _3509_/X _3511_/X _3245_/X vssd1 vssd1 vccd1 vccd1 _6125_/D sky130_fd_sc_hd__o21a_1
X_3443_ _3867_/A _3434_/Y _3424_/X _3821_/A vssd1 vssd1 vccd1 vccd1 _3443_/X sky130_fd_sc_hd__a22o_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4687__A1 _5884_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_51_wb_clk_i_A clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3374_ _3374_/A _4205_/A vssd1 vssd1 vccd1 vccd1 _3391_/B sky130_fd_sc_hd__nand2_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5113_ _5966_/Q _5116_/B vssd1 vssd1 vccd1 vccd1 _5113_/X sky130_fd_sc_hd__or2_1
XFILLER_84_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6093_ _6115_/CLK _6093_/D vssd1 vssd1 vccd1 vccd1 _6093_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _3417_/Y _3219_/X _5042_/X _5043_/X vssd1 vssd1 vccd1 vccd1 _5946_/D sky130_fd_sc_hd__o211a_1
XFILLER_53_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5946_ _5988_/CLK _5946_/D vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dfxtp_1
X_5877_ _6024_/CLK _5877_/D vssd1 vssd1 vccd1 vccd1 _5877_/Q sky130_fd_sc_hd__dfxtp_1
X_4828_ _5898_/Q _4807_/X _4826_/X _4827_/X vssd1 vssd1 vccd1 vccd1 _5898_/D sky130_fd_sc_hd__a22o_1
XFILLER_33_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4759_ _5704_/Q _5681_/Q _4797_/S vssd1 vssd1 vccd1 vccd1 _4759_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_12_wb_clk_i _5813_/CLK vssd1 vssd1 vccd1 vccd1 _5808_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_68_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5563__C1 _5556_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3634__A _3668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3090_ _3375_/B vssd1 vssd1 vccd1 vccd1 _3411_/B sky130_fd_sc_hd__buf_2
XANTENNA__3892__A2 _3287_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3992_ _3992_/A vssd1 vssd1 vccd1 vccd1 _5734_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5800_ _5959_/CLK _5800_/D vssd1 vssd1 vccd1 vccd1 _5800_/Q sky130_fd_sc_hd__dfxtp_1
X_5731_ _5808_/CLK _5731_/D vssd1 vssd1 vccd1 vccd1 _5731_/Q sky130_fd_sc_hd__dfxtp_1
X_2943_ _5285_/A _3407_/A vssd1 vssd1 vccd1 vccd1 _3003_/A sky130_fd_sc_hd__nor2_1
XFILLER_22_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2874_ _3044_/D _2950_/A _2950_/B _3312_/B vssd1 vssd1 vccd1 vccd1 _4281_/C sky130_fd_sc_hd__or4b_1
XFILLER_30_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5662_ _6109_/CLK _5662_/D vssd1 vssd1 vccd1 vccd1 _5662_/Q sky130_fd_sc_hd__dfxtp_1
X_5593_ _5393_/X _5580_/X _5592_/X _5586_/X vssd1 vssd1 vccd1 vccd1 _6101_/D sky130_fd_sc_hd__o211a_1
X_4613_ _6114_/Q _4612_/X _5624_/A vssd1 vssd1 vccd1 vccd1 _4613_/X sky130_fd_sc_hd__mux2_1
X_4544_ _4549_/A _4544_/B vssd1 vssd1 vccd1 vccd1 _5868_/D sky130_fd_sc_hd__nor2_1
Xuser_proj_example_280 vssd1 vssd1 vccd1 vccd1 io_out[28] user_proj_example_280/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_89_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4475_ _3466_/A _4469_/X _4475_/S vssd1 vssd1 vccd1 vccd1 _4476_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3426_ _5285_/A _5323_/B vssd1 vssd1 vccd1 vccd1 _5320_/A sky130_fd_sc_hd__nor2_1
X_3357_ _4321_/S vssd1 vssd1 vccd1 vccd1 _3357_/X sky130_fd_sc_hd__clkbuf_2
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6076_ _6077_/CLK _6076_/D vssd1 vssd1 vccd1 vccd1 _6076_/Q sky130_fd_sc_hd__dfxtp_1
X_3288_ _3321_/A _3322_/A _3288_/C vssd1 vssd1 vccd1 vccd1 _4470_/C sky130_fd_sc_hd__and3_1
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5027_ _5940_/Q _5030_/C vssd1 vssd1 vccd1 vccd1 _5029_/A sky130_fd_sc_hd__and2_1
XFILLER_45_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5929_ _5929_/CLK _5929_/D vssd1 vssd1 vccd1 vccd1 _5929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input22_A la_data_in[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3629__A _3632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_294 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3562__B2 _3255_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3364__A _5258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4260_ _3438_/A _3322_/X _3440_/C _4466_/B vssd1 vssd1 vccd1 vccd1 _4260_/X sky130_fd_sc_hd__a31o_1
XFILLER_79_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3211_ _6018_/Q _3208_/Y _5012_/A _6017_/Q _3210_/Y vssd1 vssd1 vccd1 vccd1 _3214_/C
+ sky130_fd_sc_hd__o221a_1
X_4191_ _5799_/Q _4190_/X _4200_/S vssd1 vssd1 vccd1 vccd1 _4192_/A sky130_fd_sc_hd__mux2_1
X_3142_ _3723_/C vssd1 vssd1 vccd1 vccd1 _5284_/A sky130_fd_sc_hd__buf_2
XFILLER_39_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3073_ _5818_/Q vssd1 vssd1 vccd1 vccd1 _3092_/C sky130_fd_sc_hd__inv_2
XFILLER_54_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3975_ _3979_/A _3975_/B vssd1 vssd1 vccd1 vccd1 _5729_/D sky130_fd_sc_hd__nor2_1
XFILLER_62_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2926_ _5323_/B _3429_/B _4438_/B vssd1 vssd1 vccd1 vccd1 _3015_/A sky130_fd_sc_hd__or3_1
XANTENNA__3250__B1 _5171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5714_ _5941_/CLK _5714_/D vssd1 vssd1 vccd1 vccd1 _5714_/Q sky130_fd_sc_hd__dfxtp_1
X_2857_ _5247_/A vssd1 vssd1 vccd1 vccd1 _2858_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5645_ _5376_/X _3576_/X _5644_/X _5638_/X vssd1 vssd1 vccd1 vccd1 _6133_/D sky130_fd_sc_hd__o211a_1
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4750__A0 _6103_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5576_ _5369_/X _5559_/A _5575_/X _5571_/X vssd1 vssd1 vccd1 vccd1 _6095_/D sky130_fd_sc_hd__o211a_1
X_4527_ _4534_/C vssd1 vssd1 vccd1 vccd1 _4527_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3274__A _3820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4458_ _4458_/A vssd1 vssd1 vccd1 vccd1 _5408_/A sky130_fd_sc_hd__buf_2
XANTENNA__3305__B2 _3117_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3305__A1 _3480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3409_ _3357_/X _3397_/X _3496_/A _3406_/Y _3408_/X vssd1 vssd1 vccd1 vccd1 _3409_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_49_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6128_ _6132_/CLK _6128_/D vssd1 vssd1 vccd1 vccd1 _6128_/Q sky130_fd_sc_hd__dfxtp_1
X_4389_ _4389_/A vssd1 vssd1 vccd1 vccd1 _5832_/D sky130_fd_sc_hd__clkbuf_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6059_ _6108_/CLK _6059_/D vssd1 vssd1 vccd1 vccd1 _6059_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4805__A1 _6036_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3440__C _3440_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_492 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_191 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3760_ _3768_/A _3760_/B vssd1 vssd1 vccd1 vccd1 _3761_/A sky130_fd_sc_hd__and2_1
XFILLER_32_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3691_ _3601_/A _5684_/Q _3697_/S vssd1 vssd1 vccd1 vccd1 _3692_/B sky130_fd_sc_hd__mux2_1
X_5430_ _6041_/Q _5439_/B vssd1 vssd1 vccd1 vccd1 _5430_/X sky130_fd_sc_hd__or2_1
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3094__A _3391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5361_ _6020_/Q _5367_/B vssd1 vssd1 vccd1 vccd1 _5361_/X sky130_fd_sc_hd__or2_1
X_5292_ _5327_/B _3424_/X _5289_/Y _5291_/X _4113_/A vssd1 vssd1 vccd1 vccd1 _5292_/X
+ sky130_fd_sc_hd__o221a_1
X_4312_ _5811_/Q _4297_/B _4311_/Y _3609_/X vssd1 vssd1 vccd1 vccd1 _5811_/D sky130_fd_sc_hd__o211a_1
XFILLER_87_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4243_ _4243_/A _4329_/B _4242_/X vssd1 vssd1 vccd1 vccd1 _4244_/A sky130_fd_sc_hd__or3b_1
XFILLER_59_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4174_ _5794_/Q _4173_/X _4184_/S vssd1 vssd1 vccd1 vccd1 _4175_/A sky130_fd_sc_hd__mux2_1
X_3125_ _5011_/A vssd1 vssd1 vccd1 vccd1 _3547_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_67_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3056_ _3857_/B vssd1 vssd1 vccd1 vccd1 _3460_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_139 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3958_ _5725_/Q _3932_/X _3957_/X vssd1 vssd1 vccd1 vccd1 _3959_/B sky130_fd_sc_hd__a21oi_1
X_2909_ _5817_/Q vssd1 vssd1 vccd1 vccd1 _2949_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_3889_ _3869_/A _3884_/X _3889_/S vssd1 vssd1 vccd1 vccd1 _3890_/A sky130_fd_sc_hd__mux2_1
X_5628_ _5342_/X _5623_/X _5626_/X _5627_/X vssd1 vssd1 vccd1 vccd1 _6113_/D sky130_fd_sc_hd__o211a_1
X_5559_ _5559_/A vssd1 vssd1 vccd1 vccd1 _5559_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3732__A _3732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5394__A _6029_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3626__B _5174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4714__B1 _4623_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5333__S _5336_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output53_A _5880_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4245__A2 _4228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5442__A1 _5366_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4930_ _6036_/Q _4924_/X _4928_/Y _4929_/X vssd1 vssd1 vccd1 vccd1 _5910_/D sky130_fd_sc_hd__o211a_1
XFILLER_52_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4861_ _5998_/Q _5990_/Q _4898_/S vssd1 vssd1 vccd1 vccd1 _4861_/X sky130_fd_sc_hd__mux2_1
X_3812_ _3810_/X _3405_/A _3812_/S vssd1 vssd1 vccd1 vccd1 _3813_/A sky130_fd_sc_hd__mux2_1
X_4792_ _6083_/Q _4834_/B vssd1 vssd1 vccd1 vccd1 _4792_/X sky130_fd_sc_hd__or2_1
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3743_ _5382_/A _5698_/Q _3753_/S vssd1 vssd1 vccd1 vccd1 _3744_/B sky130_fd_sc_hd__mux2_1
XFILLER_9_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3674_ _3674_/A vssd1 vssd1 vccd1 vccd1 _5679_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3796__D_N _3564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5413_ _6035_/Q _5417_/B vssd1 vssd1 vccd1 vccd1 _5413_/X sky130_fd_sc_hd__or2_1
X_5344_ _5348_/A vssd1 vssd1 vccd1 vccd1 _5624_/B sky130_fd_sc_hd__clkbuf_2
X_5275_ _5277_/B _5266_/X _5274_/X _5169_/X vssd1 vssd1 vccd1 vccd1 _6007_/D sky130_fd_sc_hd__o211a_1
X_4226_ _4283_/C _3845_/D _4452_/S _5255_/B _4225_/Y vssd1 vssd1 vccd1 vccd1 _4227_/C
+ sky130_fd_sc_hd__o2111a_1
XFILLER_68_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4157_ _5789_/Q _4156_/X _4167_/S vssd1 vssd1 vccd1 vccd1 _4158_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3108_ _4447_/A vssd1 vssd1 vccd1 vccd1 _5234_/A sky130_fd_sc_hd__buf_2
XFILLER_55_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4088_ _4088_/A vssd1 vssd1 vccd1 vccd1 _5769_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5479__A _6059_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5433__A1 _5353_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3039_ _3049_/A _5721_/Q vssd1 vssd1 vccd1 vccd1 _3040_/B sky130_fd_sc_hd__nand2_1
XFILLER_15_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_37_wb_clk_i clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5959_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_62_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_proj_example_109 vssd1 vssd1 vccd1 vccd1 user_proj_example_109/HI io_oeb[27]
+ sky130_fd_sc_hd__conb_1
XFILLER_7_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_451 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput14 la_data_in[40] vssd1 vssd1 vccd1 vccd1 _5376_/A sky130_fd_sc_hd__clkbuf_1
Xinput25 la_data_in[50] vssd1 vssd1 vccd1 vccd1 _3601_/A sky130_fd_sc_hd__clkbuf_1
Xinput36 la_data_in[60] vssd1 vssd1 vccd1 vccd1 _5065_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput47 wbs_stb_i vssd1 vssd1 vccd1 vccd1 _3570_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_10_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_41_wb_clk_i_A clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3390_ _3424_/B _3407_/B vssd1 vssd1 vccd1 vccd1 _3390_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__3910__A1 _5962_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5060_ _5949_/Q _5066_/B vssd1 vssd1 vccd1 vccd1 _5060_/X sky130_fd_sc_hd__or2_1
X_4011_ _4187_/A vssd1 vssd1 vccd1 vccd1 _4028_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5962_ _6064_/CLK _5962_/D vssd1 vssd1 vccd1 vccd1 _5962_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_37_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4913_ _5907_/Q _4623_/X _4911_/X _4912_/X vssd1 vssd1 vccd1 vccd1 _5907_/D sky130_fd_sc_hd__a22o_1
XANTENNA__5179__A0 _5056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5893_ _6085_/CLK _5893_/D vssd1 vssd1 vccd1 vccd1 _5893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4844_ _4819_/X _4841_/X _4843_/X _4824_/X vssd1 vssd1 vccd1 vccd1 _4844_/X sky130_fd_sc_hd__o211a_1
X_4775_ _6057_/Q _4757_/X _4767_/X _4774_/X vssd1 vssd1 vccd1 vccd1 _4775_/X sky130_fd_sc_hd__a211o_1
XANTENNA__3547__A _3547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3726_ _3732_/A _3726_/B vssd1 vssd1 vccd1 vccd1 _3727_/A sky130_fd_sc_hd__and2_1
X_3657_ _3666_/A _3657_/B vssd1 vssd1 vccd1 vccd1 _3658_/A sky130_fd_sc_hd__and2_1
X_3588_ _5046_/A _3588_/B _5046_/B vssd1 vssd1 vccd1 vccd1 _3765_/A sky130_fd_sc_hd__and3_2
X_5327_ _5327_/A _5327_/B vssd1 vssd1 vccd1 vccd1 _5327_/X sky130_fd_sc_hd__or2_1
XFILLER_0_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5258_ _5258_/A _5258_/B vssd1 vssd1 vccd1 vccd1 _5258_/Y sky130_fd_sc_hd__nor2_1
XFILLER_57_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4209_ _4209_/A vssd1 vssd1 vccd1 vccd1 _5804_/D sky130_fd_sc_hd__clkbuf_1
X_5189_ _5065_/A _5993_/Q _5189_/S vssd1 vssd1 vccd1 vccd1 _5190_/B sky130_fd_sc_hd__mux2_1
XFILLER_28_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3353__C1 _4458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4288__A _4288_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5645__A1 _5376_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_8_wb_clk_i_A _5813_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2890_ _3159_/B vssd1 vssd1 vccd1 vccd1 _3837_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_63_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4560_ _3556_/A _4529_/B _4559_/X _4460_/X vssd1 vssd1 vccd1 vccd1 _5872_/D sky130_fd_sc_hd__o211a_1
XFILLER_8_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4491_ _4562_/B _4490_/Y _4489_/B _5858_/Q vssd1 vssd1 vccd1 vccd1 _4491_/X sky130_fd_sc_hd__a211o_1
X_3511_ _3269_/X _5249_/A _5269_/A _3509_/A vssd1 vssd1 vccd1 vccd1 _3511_/X sky130_fd_sc_hd__a22o_1
X_3442_ _5247_/B vssd1 vssd1 vccd1 vccd1 _3867_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5333__A0 _6066_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3373_ _3373_/A _3373_/B vssd1 vssd1 vccd1 vccd1 _4205_/A sky130_fd_sc_hd__nand2_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3895__A0 _6112_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5112_ _5059_/X _5104_/X _5111_/X _5098_/X vssd1 vssd1 vccd1 vccd1 _5965_/D sky130_fd_sc_hd__o211a_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5636__A1 _5363_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6092_ _6115_/CLK _6092_/D vssd1 vssd1 vccd1 vccd1 _6092_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5043_ _5067_/A vssd1 vssd1 vccd1 vccd1 _5043_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__3647__A0 _5369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5945_ _5945_/CLK _5945_/D vssd1 vssd1 vccd1 vccd1 _5945_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5876_ _5945_/CLK _5876_/D vssd1 vssd1 vccd1 vccd1 _5876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4827_ _6038_/Q _4803_/X _4804_/X vssd1 vssd1 vccd1 vccd1 _4827_/X sky130_fd_sc_hd__o21a_1
XFILLER_21_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4758_ _4860_/A vssd1 vssd1 vccd1 vccd1 _4797_/S sky130_fd_sc_hd__clkbuf_2
X_3709_ _3709_/A vssd1 vssd1 vccd1 vccd1 _5689_/D sky130_fd_sc_hd__clkbuf_1
X_4689_ _6133_/Q _4688_/X _4719_/S vssd1 vssd1 vccd1 vccd1 _4689_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5492__A _5535_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3638__A0 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_52_wb_clk_i clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6027_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_16_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3810__A0 _6058_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3892__A3 _3466_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3650__A _3668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3991_ _3994_/A _3991_/B vssd1 vssd1 vccd1 vccd1 _3992_/A sky130_fd_sc_hd__and2_1
XFILLER_74_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5730_ _5736_/CLK _5730_/D vssd1 vssd1 vccd1 vccd1 _5730_/Q sky130_fd_sc_hd__dfxtp_1
X_2942_ _2942_/A vssd1 vssd1 vccd1 vccd1 _3407_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2873_ _5816_/Q vssd1 vssd1 vccd1 vccd1 _3312_/B sky130_fd_sc_hd__clkbuf_1
X_5661_ _6108_/CLK _5661_/D vssd1 vssd1 vccd1 vccd1 _5661_/Q sky130_fd_sc_hd__dfxtp_1
X_5592_ _6101_/Q _5592_/B vssd1 vssd1 vccd1 vccd1 _5592_/X sky130_fd_sc_hd__or2_1
X_4612_ _5690_/Q _5667_/Q _4645_/S vssd1 vssd1 vccd1 vccd1 _4612_/X sky130_fd_sc_hd__mux2_1
X_4543_ _4545_/B _4545_/C vssd1 vssd1 vccd1 vccd1 _4544_/B sky130_fd_sc_hd__xnor2_1
Xuser_proj_example_281 vssd1 vssd1 vccd1 vccd1 io_out[29] user_proj_example_281/LO
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_270 vssd1 vssd1 vccd1 vccd1 io_out[18] user_proj_example_270/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA__5306__B1 _4041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4474_ _4555_/B _4555_/C _4474_/C _4556_/C vssd1 vssd1 vccd1 vccd1 _4475_/S sky130_fd_sc_hd__and4bb_1
X_3425_ _3275_/X _3423_/X _3424_/X _3360_/X vssd1 vssd1 vccd1 vccd1 _3425_/X sky130_fd_sc_hd__a2bb2o_1
XANTENNA__3868__B1 _5761_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3356_ _3354_/X _3355_/X _4322_/A vssd1 vssd1 vccd1 vccd1 _3356_/X sky130_fd_sc_hd__a21o_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3287_ _4470_/A vssd1 vssd1 vccd1 vccd1 _3287_/X sky130_fd_sc_hd__buf_2
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6075_ _6135_/CLK _6075_/D vssd1 vssd1 vccd1 vccd1 _6075_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5026_ _5026_/A vssd1 vssd1 vccd1 vccd1 _5939_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_535 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4045__A0 _6099_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5928_ _5945_/CLK _5928_/D vssd1 vssd1 vccd1 vccd1 _5928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5859_ _5874_/CLK _5859_/D vssd1 vssd1 vccd1 vccd1 _5859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4566__A _5188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input15_A la_data_in[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5397__A _6030_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4339__A1 _3275_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5336__S _5336_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4448__A1_N _3897_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3210_ _6019_/Q _5938_/Q vssd1 vssd1 vccd1 vccd1 _3210_/Y sky130_fd_sc_hd__xnor2_1
X_4190_ _5949_/Q _5798_/Q _4196_/S vssd1 vssd1 vccd1 vccd1 _4190_/X sky130_fd_sc_hd__mux2_1
X_3141_ _3408_/B vssd1 vssd1 vccd1 vccd1 _3723_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_39_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3380__A _5234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3072_ _3824_/A _5818_/Q vssd1 vssd1 vccd1 vccd1 _3349_/C sky130_fd_sc_hd__nor2_1
XFILLER_54_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3974_ _5729_/Q _3932_/X _3973_/X vssd1 vssd1 vccd1 vccd1 _3975_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__5100__A _5962_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2925_ _2959_/C _3465_/B _3044_/D _3465_/C vssd1 vssd1 vccd1 vccd1 _4438_/B sky130_fd_sc_hd__nand4b_4
X_5713_ _5892_/CLK _5713_/D vssd1 vssd1 vccd1 vccd1 _5713_/Q sky130_fd_sc_hd__dfxtp_2
X_2856_ _4281_/A vssd1 vssd1 vccd1 vccd1 _5247_/A sky130_fd_sc_hd__clkbuf_2
X_5644_ _6133_/Q _5648_/B vssd1 vssd1 vccd1 vccd1 _5644_/X sky130_fd_sc_hd__or2_1
X_5575_ _6095_/Q _5577_/B vssd1 vssd1 vccd1 vccd1 _5575_/X sky130_fd_sc_hd__or2_1
X_4526_ _5742_/Q _5738_/Q _5737_/Q _4500_/Y vssd1 vssd1 vccd1 vccd1 _4534_/C sky130_fd_sc_hd__o31a_1
X_4457_ _5248_/A _5249_/A _3505_/C _3390_/Y _4567_/A vssd1 vssd1 vccd1 vccd1 _4457_/X
+ sky130_fd_sc_hd__a41o_1
X_3408_ _3513_/B _3408_/B _4366_/A vssd1 vssd1 vccd1 vccd1 _3408_/X sky130_fd_sc_hd__or3b_1
XANTENNA__3305__A2 _3459_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6127_ _6131_/CLK _6127_/D vssd1 vssd1 vccd1 vccd1 _6127_/Q sky130_fd_sc_hd__dfxtp_1
X_4388_ _5832_/Q _4387_/X _4391_/S vssd1 vssd1 vccd1 vccd1 _4389_/A sky130_fd_sc_hd__mux2_1
XANTENNA_input7_A la_data_in[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3339_ _3853_/A _3493_/A vssd1 vssd1 vccd1 vccd1 _4293_/A sky130_fd_sc_hd__xor2_2
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6058_ _6108_/CLK _6058_/D vssd1 vssd1 vccd1 vccd1 _6058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5009_ _5935_/Q _5008_/A _4995_/B vssd1 vssd1 vccd1 vccd1 _5009_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_26_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3690_ _3690_/A vssd1 vssd1 vccd1 vccd1 _5683_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3375__A _3553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5360_ input8/X vssd1 vssd1 vccd1 vccd1 _5360_/X sky130_fd_sc_hd__clkbuf_2
X_5291_ _5323_/A _5246_/B _5290_/X _3867_/A vssd1 vssd1 vccd1 vccd1 _5291_/X sky130_fd_sc_hd__o211a_1
X_4311_ _4307_/Y _4309_/X _4310_/X vssd1 vssd1 vccd1 vccd1 _4311_/Y sky130_fd_sc_hd__o21ai_1
X_4242_ _4294_/A _4294_/B _4242_/C vssd1 vssd1 vccd1 vccd1 _4242_/X sky130_fd_sc_hd__and3_1
XFILLER_4_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5590__A _6100_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4173_ _5662_/Q _5793_/Q _4179_/S vssd1 vssd1 vccd1 vccd1 _4173_/X sky130_fd_sc_hd__mux2_1
X_3124_ _3423_/B vssd1 vssd1 vccd1 vccd1 _5011_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_67_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3055_ _5241_/A _3841_/B _3037_/B _3451_/D vssd1 vssd1 vccd1 vccd1 _3055_/X sky130_fd_sc_hd__o31a_1
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3471__A1 _5279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3471__B2 _3854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_482 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3957_ _5724_/Q _3941_/X _3953_/X _3956_/Y vssd1 vssd1 vccd1 vccd1 _3957_/X sky130_fd_sc_hd__o211a_1
XFILLER_23_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2908_ _2950_/A vssd1 vssd1 vccd1 vccd1 _3322_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_50_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3888_ _3888_/A _5236_/B vssd1 vssd1 vccd1 vccd1 _3889_/S sky130_fd_sc_hd__nor2_1
XFILLER_31_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2839_ _6012_/Q vssd1 vssd1 vccd1 vccd1 _5327_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5627_ _5638_/A vssd1 vssd1 vccd1 vccd1 _5627_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3526__A2 _4331_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5558_ _5601_/B _5622_/B vssd1 vssd1 vccd1 vccd1 _5559_/A sky130_fd_sc_hd__or2_1
X_4509_ _4518_/D _4506_/B _4518_/C vssd1 vssd1 vccd1 vccd1 _4512_/B sky130_fd_sc_hd__a21oi_1
XFILLER_2_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5489_ _3614_/X _5470_/A _5487_/X _5488_/X vssd1 vssd1 vccd1 vccd1 _6063_/D sky130_fd_sc_hd__o211a_1
XFILLER_76_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_31_wb_clk_i_A _5836_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4714__A1 _5387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_7_wb_clk_i _5813_/CLK vssd1 vssd1 vccd1 vccd1 _5796_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_1_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5288__C _5301_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4860_ _4860_/A vssd1 vssd1 vccd1 vccd1 _4898_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_32_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3811_ _4383_/A _3379_/A _3525_/A vssd1 vssd1 vccd1 vccd1 _3812_/S sky130_fd_sc_hd__o21ai_2
XFILLER_20_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4791_ _4842_/A vssd1 vssd1 vccd1 vccd1 _4834_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_20_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5585__A _6098_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3742_ _3742_/A vssd1 vssd1 vccd1 vccd1 _5697_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3673_ _3684_/A _3673_/B vssd1 vssd1 vccd1 vccd1 _3674_/A sky130_fd_sc_hd__and2_1
X_5412_ _3598_/X _5404_/X _5411_/X _5409_/X vssd1 vssd1 vccd1 vccd1 _6034_/D sky130_fd_sc_hd__o211a_1
X_5343_ _5343_/A _5343_/B vssd1 vssd1 vccd1 vccd1 _5348_/A sky130_fd_sc_hd__nand2_1
X_5274_ _5274_/A _5274_/B _5294_/S vssd1 vssd1 vccd1 vccd1 _5274_/X sky130_fd_sc_hd__or3b_1
XFILLER_68_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4225_ _3834_/B _4220_/Y _4224_/X vssd1 vssd1 vccd1 vccd1 _4225_/Y sky130_fd_sc_hd__a21oi_1
X_4156_ _5656_/Q _5788_/Q _4162_/S vssd1 vssd1 vccd1 vccd1 _4156_/X sky130_fd_sc_hd__mux2_1
X_3107_ _3814_/B vssd1 vssd1 vccd1 vccd1 _4447_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4087_ _5769_/Q _4086_/X _4097_/S vssd1 vssd1 vccd1 vccd1 _4088_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4664__A _4716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3038_ _3038_/A _5721_/Q vssd1 vssd1 vccd1 vccd1 _3463_/B sky130_fd_sc_hd__or2_1
XFILLER_23_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4989_ _4989_/A vssd1 vssd1 vccd1 vccd1 _5928_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3462__B _3480_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4293__B _4327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput15 la_data_in[41] vssd1 vssd1 vccd1 vccd1 _5382_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput26 la_data_in[51] vssd1 vssd1 vccd1 vccd1 _3604_/A sky130_fd_sc_hd__clkbuf_1
Xinput37 la_data_in[61] vssd1 vssd1 vccd1 vccd1 _5069_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput48 wbs_we_i vssd1 vssd1 vccd1 vccd1 _5046_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_6_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4699__A0 _6098_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3910__A2 _3061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4010_ _4010_/A _4473_/B vssd1 vssd1 vccd1 vccd1 _4187_/A sky130_fd_sc_hd__nor2_1
XFILLER_37_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5961_ _6064_/CLK _5961_/D vssd1 vssd1 vccd1 vccd1 _5961_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4912_ _5985_/Q _5379_/B _4607_/A vssd1 vssd1 vccd1 vccd1 _4912_/X sky130_fd_sc_hd__o21a_1
X_5892_ _5892_/CLK _5892_/D vssd1 vssd1 vccd1 vccd1 _5892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4843_ _6088_/Q _4885_/B vssd1 vssd1 vccd1 vccd1 _4843_/X sky130_fd_sc_hd__or2_1
XANTENNA__4926__A1 _6035_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4774_ _4768_/X _4771_/X _4772_/X _4773_/X vssd1 vssd1 vccd1 vccd1 _4774_/X sky130_fd_sc_hd__o211a_1
X_3725_ input9/X _5693_/Q _3735_/S vssd1 vssd1 vccd1 vccd1 _3726_/B sky130_fd_sc_hd__mux2_1
X_3656_ _5376_/A _5674_/Q _3669_/S vssd1 vssd1 vccd1 vccd1 _3657_/B sky130_fd_sc_hd__mux2_1
X_3587_ _3587_/A vssd1 vssd1 vccd1 vccd1 _3587_/X sky130_fd_sc_hd__clkbuf_2
X_5326_ _5244_/B _5320_/Y _5322_/X _5325_/X vssd1 vssd1 vccd1 vccd1 _5326_/X sky130_fd_sc_hd__a31o_1
XANTENNA_clkbuf_3_6__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5257_ _5257_/A _5257_/B vssd1 vssd1 vccd1 vccd1 _5257_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4457__A3 _3505_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4208_ _4524_/A _4208_/B vssd1 vssd1 vccd1 vccd1 _4209_/A sky130_fd_sc_hd__and2_1
XFILLER_87_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5188_ _5188_/A vssd1 vssd1 vccd1 vccd1 _5204_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4139_ _6134_/Q _5783_/Q _4145_/S vssd1 vssd1 vccd1 vccd1 _4139_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3738__A _3738_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input45_A wbs_sel_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3367__B _3891_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3510_ _3424_/B _3407_/B _6125_/Q vssd1 vssd1 vccd1 vccd1 _5269_/A sky130_fd_sc_hd__o21a_1
X_4490_ _5743_/Q vssd1 vssd1 vccd1 vccd1 _4490_/Y sky130_fd_sc_hd__inv_2
X_3441_ _3326_/A _3429_/X _3031_/Y _2936_/A _3440_/X vssd1 vssd1 vccd1 vccd1 _3441_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_6_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3372_ _3935_/C _6125_/Q _3469_/A vssd1 vssd1 vccd1 vccd1 _3372_/X sky130_fd_sc_hd__o21a_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5111_ _5965_/Q _5116_/B vssd1 vssd1 vccd1 vccd1 _5111_/X sky130_fd_sc_hd__or2_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6091_ _6091_/CLK _6091_/D vssd1 vssd1 vccd1 vccd1 _6091_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5042_ _5854_/Q _3218_/X _3135_/A vssd1 vssd1 vccd1 vccd1 _5042_/X sky130_fd_sc_hd__a21o_1
XFILLER_84_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5103__A _5535_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5944_ _5944_/CLK _5944_/D vssd1 vssd1 vccd1 vccd1 _5944_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5875_ _5945_/CLK _5875_/D vssd1 vssd1 vccd1 vccd1 _5875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4826_ _6062_/Q _4808_/X _4818_/X _4825_/X vssd1 vssd1 vccd1 vccd1 _4826_/X sky130_fd_sc_hd__a211o_1
X_4757_ _4859_/A vssd1 vssd1 vccd1 vccd1 _4757_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__5572__A1 _5363_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3708_ _3732_/A _3708_/B vssd1 vssd1 vccd1 vccd1 _3709_/A sky130_fd_sc_hd__and2_1
X_4688_ _5697_/Q _5674_/Q _4697_/S vssd1 vssd1 vccd1 vccd1 _4688_/X sky130_fd_sc_hd__mux2_1
X_3639_ _3648_/A _3639_/B vssd1 vssd1 vccd1 vccd1 _3640_/A sky130_fd_sc_hd__and2_1
X_5309_ _5309_/A vssd1 vssd1 vccd1 vccd1 _5315_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_396 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_21_wb_clk_i clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6121_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4599__C1 _5469_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4063__S _4063_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3169__A3 _3484_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5563__A1 _5342_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3990_ _5734_/Q _3964_/X _3953_/A _5733_/Q vssd1 vssd1 vccd1 vccd1 _3991_/B sky130_fd_sc_hd__a22o_1
XFILLER_62_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2941_ _2941_/A vssd1 vssd1 vccd1 vccd1 _5285_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_15_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3378__A _6121_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5660_ _6108_/CLK _5660_/D vssd1 vssd1 vccd1 vccd1 _5660_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2872_ _5817_/Q vssd1 vssd1 vccd1 vccd1 _2950_/B sky130_fd_sc_hd__clkbuf_1
X_4611_ _4717_/A vssd1 vssd1 vccd1 vccd1 _4611_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5554__A1 _3614_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5591_ _5389_/X _5580_/X _5590_/X _5586_/X vssd1 vssd1 vccd1 vccd1 _6100_/D sky130_fd_sc_hd__o211a_1
X_4542_ _4549_/A _4542_/B _4545_/C vssd1 vssd1 vccd1 vccd1 _5867_/D sky130_fd_sc_hd__nor3_1
Xuser_proj_example_282 vssd1 vssd1 vccd1 vccd1 io_out[30] user_proj_example_282/LO
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_271 vssd1 vssd1 vccd1 vccd1 io_out[19] user_proj_example_271/LO
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_260 vssd1 vssd1 vccd1 vccd1 io_out[8] user_proj_example_260/LO
+ sky130_fd_sc_hd__conb_1
X_4473_ _5254_/B _4473_/B _3901_/Y vssd1 vssd1 vccd1 vccd1 _4556_/C sky130_fd_sc_hd__nor3b_1
XFILLER_7_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3424_ _3429_/B _3424_/B vssd1 vssd1 vccd1 vccd1 _3424_/X sky130_fd_sc_hd__or2_1
XANTENNA__4002__A _4002_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3868__A1 _3869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3355_ _6130_/Q _5818_/Q _5715_/Q _4235_/C vssd1 vssd1 vccd1 vccd1 _3355_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3841__A _3841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3286_ _5719_/Q vssd1 vssd1 vccd1 vccd1 _4470_/A sky130_fd_sc_hd__clkbuf_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6074_ _6080_/CLK _6074_/D vssd1 vssd1 vccd1 vccd1 _6074_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5025_ _5030_/C _5025_/B _5025_/C vssd1 vssd1 vccd1 vccd1 _5026_/A sky130_fd_sc_hd__and3b_1
XFILLER_26_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5927_ _5944_/CLK _5927_/D vssd1 vssd1 vccd1 vccd1 _5927_/Q sky130_fd_sc_hd__dfxtp_1
X_5858_ _6131_/CLK _5858_/D vssd1 vssd1 vccd1 vccd1 _5858_/Q sky130_fd_sc_hd__dfxtp_1
X_4809_ _4860_/A vssd1 vssd1 vccd1 vccd1 _4848_/S sky130_fd_sc_hd__clkbuf_2
X_5789_ _6115_/CLK _5789_/D vssd1 vssd1 vccd1 vccd1 _5789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_403 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4284__A1 _3480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3795__B1 _3411_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4757__A _4859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3140_ _3411_/B vssd1 vssd1 vccd1 vccd1 _3408_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_67_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3071_ _3071_/A vssd1 vssd1 vccd1 vccd1 _3274_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5588__A _6099_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3973_ _5728_/Q _3941_/X _3953_/X _3972_/Y vssd1 vssd1 vccd1 vccd1 _3973_/X sky130_fd_sc_hd__o211a_1
XFILLER_62_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5712_ _6087_/CLK _5712_/D vssd1 vssd1 vccd1 vccd1 _5712_/Q sky130_fd_sc_hd__dfxtp_1
X_2924_ _3312_/D vssd1 vssd1 vccd1 vccd1 _3465_/C sky130_fd_sc_hd__clkbuf_2
X_2855_ _3845_/A vssd1 vssd1 vccd1 vccd1 _4281_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5527__A1 _5393_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5643_ _5373_/X _5623_/A _5642_/X _5638_/X vssd1 vssd1 vccd1 vccd1 _6120_/D sky130_fd_sc_hd__o211a_1
XANTENNA__3836__A _3836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5574_ _5366_/X _5559_/A _5573_/X _5571_/X vssd1 vssd1 vccd1 vccd1 _6094_/D sky130_fd_sc_hd__o211a_1
X_4525_ _4525_/A vssd1 vssd1 vccd1 vccd1 _5864_/D sky130_fd_sc_hd__clkbuf_1
X_4456_ _3469_/A _5249_/A _5248_/A _3269_/X vssd1 vssd1 vccd1 vccd1 _4456_/X sky130_fd_sc_hd__a211o_1
X_3407_ _3407_/A _3407_/B vssd1 vssd1 vccd1 vccd1 _3513_/B sky130_fd_sc_hd__or2_2
X_4387_ _6054_/Q _5831_/Q _4396_/S vssd1 vssd1 vccd1 vccd1 _4387_/X sky130_fd_sc_hd__mux2_1
X_6126_ _6132_/CLK _6126_/D vssd1 vssd1 vccd1 vccd1 _6126_/Q sky130_fd_sc_hd__dfxtp_1
X_3338_ _5714_/Q vssd1 vssd1 vccd1 vccd1 _3493_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_58_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3571__A _5667_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_458 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3269_ _4206_/A vssd1 vssd1 vccd1 vccd1 _3269_/X sky130_fd_sc_hd__clkbuf_2
X_6057_ _6108_/CLK _6057_/D vssd1 vssd1 vccd1 vccd1 _6057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5008_ _5008_/A _5008_/B vssd1 vssd1 vccd1 vccd1 _5934_/D sky130_fd_sc_hd__nor2_1
XANTENNA__5498__A _6066_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4974__C1 _5284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_21_wb_clk_i_A clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_39_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4009__A1 _5284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_60_wb_clk_i_A clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_9_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3375__B _3375_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5290_ _5297_/C _5280_/A _5297_/B vssd1 vssd1 vccd1 vccd1 _5290_/X sky130_fd_sc_hd__a21o_1
X_4310_ _3494_/Y _4294_/D _4309_/X _4297_/B vssd1 vssd1 vccd1 vccd1 _4310_/X sky130_fd_sc_hd__o31a_1
X_4241_ _4241_/A _4293_/A vssd1 vssd1 vccd1 vccd1 _4242_/C sky130_fd_sc_hd__or2_1
XFILLER_4_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3391__A _3391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4172_ _4172_/A vssd1 vssd1 vccd1 vccd1 _5793_/D sky130_fd_sc_hd__clkbuf_1
X_3123_ _3508_/B _3100_/Y _3122_/X vssd1 vssd1 vccd1 vccd1 _3123_/Y sky130_fd_sc_hd__a21oi_1
X_3054_ _3054_/A _3116_/A vssd1 vssd1 vccd1 vccd1 _3451_/D sky130_fd_sc_hd__or2_1
XFILLER_67_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3956_ _5724_/Q _3983_/B vssd1 vssd1 vccd1 vccd1 _3956_/Y sky130_fd_sc_hd__nand2_1
XFILLER_50_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2907_ _4255_/A _3315_/B vssd1 vssd1 vccd1 vccd1 _4210_/B sky130_fd_sc_hd__or2_1
X_3887_ _3459_/D _3821_/X _3886_/Y vssd1 vssd1 vccd1 vccd1 _5236_/B sky130_fd_sc_hd__a21o_1
X_5626_ _6113_/Q _5635_/B vssd1 vssd1 vccd1 vccd1 _5626_/X sky130_fd_sc_hd__or2_1
X_2838_ _5277_/A vssd1 vssd1 vccd1 vccd1 _5281_/A sky130_fd_sc_hd__clkbuf_1
X_5557_ _3617_/X _5536_/A _5555_/X _5556_/X vssd1 vssd1 vccd1 vccd1 _6088_/D sky130_fd_sc_hd__o211a_1
X_4508_ _5861_/Q vssd1 vssd1 vccd1 vccd1 _4518_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5488_ _5529_/A vssd1 vssd1 vccd1 vccd1 _5488_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_78_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4439_ _3052_/A _2917_/A _3873_/D _6005_/Q _3874_/A vssd1 vssd1 vccd1 vccd1 _4439_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_58_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6109_ _6109_/CLK _6109_/D vssd1 vssd1 vccd1 vccd1 _6109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3476__A _5279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3922__A0 _3037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4478__A1 _5336_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_442 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3810_ _6058_/Q _3809_/X _5278_/A vssd1 vssd1 vccd1 vccd1 _3810_/X sky130_fd_sc_hd__mux2_1
X_4790_ _6107_/Q _4789_/X _4822_/S vssd1 vssd1 vccd1 vccd1 _4790_/X sky130_fd_sc_hd__mux2_1
X_3741_ _3750_/A _3741_/B vssd1 vssd1 vccd1 vccd1 _3742_/A sky130_fd_sc_hd__and2_1
XFILLER_20_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3672_ _5396_/A _5679_/Q _3678_/S vssd1 vssd1 vccd1 vccd1 _3673_/B sky130_fd_sc_hd__mux2_1
X_5411_ _6034_/Q _5417_/B vssd1 vssd1 vccd1 vccd1 _5411_/X sky130_fd_sc_hd__or2_1
X_5342_ input5/X vssd1 vssd1 vccd1 vccd1 _5342_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_87_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5273_ _5301_/C _5245_/B _5271_/Y _5272_/X _4041_/S vssd1 vssd1 vccd1 vccd1 _5274_/B
+ sky130_fd_sc_hd__o311a_1
XANTENNA__4469__A1 _5954_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4224_ _4447_/C _4447_/D _3849_/C vssd1 vssd1 vccd1 vccd1 _4224_/X sky130_fd_sc_hd__o21a_1
X_4155_ _4155_/A vssd1 vssd1 vccd1 vccd1 _5788_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3106_ _4231_/A vssd1 vssd1 vccd1 vccd1 _4554_/S sky130_fd_sc_hd__clkbuf_4
X_4086_ _5955_/Q _3287_/X _4092_/S vssd1 vssd1 vccd1 vccd1 _4086_/X sky130_fd_sc_hd__mux2_1
X_3037_ _3037_/A _3037_/B vssd1 vssd1 vccd1 vccd1 _3037_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4156__S _4162_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4988_ _4993_/C _4995_/B _4988_/C vssd1 vssd1 vccd1 vccd1 _4989_/A sky130_fd_sc_hd__and3b_1
XFILLER_51_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3939_ _3939_/A _3930_/A vssd1 vssd1 vccd1 vccd1 _3940_/B sky130_fd_sc_hd__or2b_1
Xclkbuf_leaf_46_wb_clk_i clkbuf_3_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6087_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_5609_ _6107_/Q _5614_/B vssd1 vssd1 vccd1 vccd1 _5609_/X sky130_fd_sc_hd__or2_1
XFILLER_3_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4855__A _4855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput16 la_data_in[42] vssd1 vssd1 vccd1 vccd1 _5386_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput27 la_data_in[52] vssd1 vssd1 vccd1 vccd1 _3607_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_6_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput38 la_data_in[62] vssd1 vssd1 vccd1 vccd1 _5072_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3145__S _5666_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5960_ _5975_/CLK _5960_/D vssd1 vssd1 vccd1 vccd1 _5960_/Q sky130_fd_sc_hd__dfxtp_1
X_5891_ _5892_/CLK _5891_/D vssd1 vssd1 vccd1 vccd1 _5891_/Q sky130_fd_sc_hd__dfxtp_1
X_4911_ _5977_/Q _4706_/A _4869_/X _4910_/X vssd1 vssd1 vccd1 vccd1 _4911_/X sky130_fd_sc_hd__a211o_1
XANTENNA__5596__A _6103_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4387__A0 _6054_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4842_ _4842_/A vssd1 vssd1 vccd1 vccd1 _4885_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4773_ _4824_/A vssd1 vssd1 vccd1 vccd1 _4773_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3724_ _3724_/A vssd1 vssd1 vccd1 vccd1 _5692_/D sky130_fd_sc_hd__clkinv_2
X_3655_ _3678_/S vssd1 vssd1 vccd1 vccd1 _3669_/S sky130_fd_sc_hd__clkbuf_2
X_3586_ _3582_/X _3576_/X _3583_/X _3585_/X vssd1 vssd1 vccd1 vccd1 _5657_/D sky130_fd_sc_hd__o211a_1
X_5325_ _5323_/X _5246_/B _5324_/X _3867_/X vssd1 vssd1 vccd1 vccd1 _5325_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5256_ _5256_/A _5256_/B _5287_/B vssd1 vssd1 vccd1 vccd1 _5257_/B sky130_fd_sc_hd__or3_1
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4207_ _4455_/A _3522_/A _5248_/B _4206_/X _5804_/Q vssd1 vssd1 vccd1 vccd1 _4208_/B
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4675__A _4855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5187_ _5187_/A vssd1 vssd1 vccd1 vccd1 _5992_/D sky130_fd_sc_hd__clkbuf_1
X_4138_ _4138_/A vssd1 vssd1 vccd1 vccd1 _5783_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4069_ _6107_/Q _5763_/Q _4075_/S vssd1 vssd1 vccd1 vccd1 _4069_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input38_A la_data_in[62] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5318__C1 _5169_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3440_ _3440_/A _3440_/B _3440_/C _3440_/D vssd1 vssd1 vccd1 vccd1 _3440_/X sky130_fd_sc_hd__and4_1
X_3371_ _6127_/Q vssd1 vssd1 vccd1 vccd1 _3935_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5110_ _5056_/X _5104_/X _5109_/X _5098_/X vssd1 vssd1 vccd1 vccd1 _5964_/D sky130_fd_sc_hd__o211a_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6090_ _6115_/CLK _6090_/D vssd1 vssd1 vccd1 vccd1 _6090_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _5945_/Q _5011_/B _3221_/X vssd1 vssd1 vccd1 vccd1 _5945_/D sky130_fd_sc_hd__o21a_1
XFILLER_84_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_92_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5943_ _5944_/CLK _5943_/D vssd1 vssd1 vccd1 vccd1 _5943_/Q sky130_fd_sc_hd__dfxtp_1
X_5874_ _5874_/CLK _5874_/D vssd1 vssd1 vccd1 vccd1 _5874_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_21_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4825_ _4819_/X _4822_/X _4823_/X _4824_/X vssd1 vssd1 vccd1 vccd1 _4825_/X sky130_fd_sc_hd__o211a_1
XANTENNA__5557__C1 _5556_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4756_ _4756_/A vssd1 vssd1 vccd1 vccd1 _4756_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3707_ _3617_/A _5689_/Q _3707_/S vssd1 vssd1 vccd1 vccd1 _3708_/B sky130_fd_sc_hd__mux2_1
X_4687_ _5884_/Q _4653_/X _4685_/X _4686_/X vssd1 vssd1 vccd1 vccd1 _5884_/D sky130_fd_sc_hd__a22o_1
X_3638_ input8/X _5669_/Q _3641_/S vssd1 vssd1 vccd1 vccd1 _3639_/B sky130_fd_sc_hd__mux2_1
X_3569_ _5624_/A vssd1 vssd1 vccd1 vccd1 _5622_/A sky130_fd_sc_hd__clkbuf_2
X_5308_ _5297_/A _5266_/X _5307_/X _5169_/X vssd1 vssd1 vccd1 vccd1 _6010_/D sky130_fd_sc_hd__o211a_1
XFILLER_68_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5239_ _5277_/C vssd1 vssd1 vccd1 vccd1 _5243_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3425__A1_N _3275_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_61_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6138_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4771__A0 _6105_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2940_ _3053_/A vssd1 vssd1 vccd1 vccd1 _3849_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_50_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2871_ _5815_/Q vssd1 vssd1 vccd1 vccd1 _2950_/A sky130_fd_sc_hd__clkbuf_1
X_4610_ _4716_/A vssd1 vssd1 vccd1 vccd1 _4610_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5590_ _6100_/Q _5592_/B vssd1 vssd1 vccd1 vccd1 _5590_/X sky130_fd_sc_hd__or2_1
X_4541_ _4541_/A _4541_/B vssd1 vssd1 vccd1 vccd1 _4545_/C sky130_fd_sc_hd__and2_1
XFILLER_7_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_proj_example_272 vssd1 vssd1 vccd1 vccd1 io_out[20] user_proj_example_272/LO
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_261 vssd1 vssd1 vccd1 vccd1 io_out[9] user_proj_example_261/LO
+ sky130_fd_sc_hd__conb_1
X_4472_ _5250_/A _3851_/C _4470_/X _4471_/Y vssd1 vssd1 vccd1 vccd1 _5254_/B sky130_fd_sc_hd__a31o_1
XFILLER_7_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xuser_proj_example_250 vssd1 vssd1 vccd1 vccd1 user_proj_example_250/HI wbs_dat_o[29]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_283 vssd1 vssd1 vccd1 vccd1 io_out[31] user_proj_example_283/LO
+ sky130_fd_sc_hd__conb_1
X_3423_ _3423_/A _3423_/B _3423_/C _3423_/D vssd1 vssd1 vccd1 vccd1 _3423_/X sky130_fd_sc_hd__or4_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3354_ _3897_/A vssd1 vssd1 vccd1 vccd1 _3354_/X sky130_fd_sc_hd__clkbuf_2
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3285_ _3350_/B vssd1 vssd1 vccd1 vccd1 _3291_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6073_ _6080_/CLK _6073_/D vssd1 vssd1 vccd1 vccd1 _6073_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5024_ _5938_/Q _5023_/C _5939_/Q vssd1 vssd1 vccd1 vccd1 _5025_/C sky130_fd_sc_hd__a21o_1
X_5926_ _5926_/CLK _5926_/D vssd1 vssd1 vccd1 vccd1 _5926_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3569__A _5624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5857_ _6121_/CLK _5857_/D vssd1 vssd1 vccd1 vccd1 _5857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_11_wb_clk_i_A _5813_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4808_ _4859_/A vssd1 vssd1 vccd1 vccd1 _4808_/X sky130_fd_sc_hd__clkbuf_2
X_5788_ _6118_/CLK _5788_/D vssd1 vssd1 vccd1 vccd1 _5788_/Q sky130_fd_sc_hd__dfxtp_1
X_4739_ _6102_/Q _4738_/X _4771_/S vssd1 vssd1 vccd1 vccd1 _4739_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4339__S _4399_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_50_wb_clk_i_A clkbuf_3_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3070_ _3266_/A vssd1 vssd1 vccd1 vccd1 _3274_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4773__A _4824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_378 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3972_ _5728_/Q _3983_/B vssd1 vssd1 vccd1 vccd1 _3972_/Y sky130_fd_sc_hd__nand2_1
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5711_ _6087_/CLK _5711_/D vssd1 vssd1 vccd1 vccd1 _5711_/Q sky130_fd_sc_hd__dfxtp_1
X_2923_ _2949_/D vssd1 vssd1 vccd1 vccd1 _3465_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_2854_ _6122_/Q vssd1 vssd1 vccd1 vccd1 _3845_/A sky130_fd_sc_hd__inv_2
X_5642_ _6120_/Q _5642_/B vssd1 vssd1 vccd1 vccd1 _5642_/X sky130_fd_sc_hd__or2_1
XANTENNA__3836__B _4288_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5573_ _6094_/Q _5577_/B vssd1 vssd1 vccd1 vccd1 _5573_/X sky130_fd_sc_hd__or2_1
X_4524_ _4524_/A _4524_/B vssd1 vssd1 vccd1 vccd1 _4525_/A sky130_fd_sc_hd__and2_1
X_4455_ _4455_/A vssd1 vssd1 vccd1 vccd1 _5248_/A sky130_fd_sc_hd__inv_2
X_3406_ _3402_/Y _3484_/B _3405_/X vssd1 vssd1 vccd1 vccd1 _3406_/Y sky130_fd_sc_hd__o21ai_4
X_4386_ _4386_/A vssd1 vssd1 vccd1 vccd1 _5831_/D sky130_fd_sc_hd__clkbuf_1
X_6125_ _6132_/CLK _6125_/D vssd1 vssd1 vccd1 vccd1 _6125_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3337_ _5856_/Q _3257_/A _3336_/X _3841_/A vssd1 vssd1 vccd1 vccd1 _3814_/C sky130_fd_sc_hd__o2bb2a_1
XANTENNA__3571__B _3794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4159__S _4162_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4266__A2 _3480_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3268_ _3800_/A vssd1 vssd1 vccd1 vccd1 _3891_/B sky130_fd_sc_hd__clkbuf_2
X_6056_ _6080_/CLK _6056_/D vssd1 vssd1 vccd1 vccd1 _6056_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3199_ _6018_/Q vssd1 vssd1 vccd1 vccd1 _5354_/A sky130_fd_sc_hd__clkinv_2
XFILLER_38_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5007_ _5934_/Q _5005_/A _4990_/X vssd1 vssd1 vccd1 vccd1 _5008_/B sky130_fd_sc_hd__o21ai_1
XFILLER_26_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5909_ _5922_/CLK _5909_/D vssd1 vssd1 vccd1 vccd1 _5909_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4858__A _4858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3481__B _3481_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input20_A la_data_in[46] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5201__B _5201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4768__A _4870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4240_ _6130_/Q _4240_/B vssd1 vssd1 vccd1 vccd1 _4294_/B sky130_fd_sc_hd__nand2_1
X_4171_ _5793_/Q _4169_/X _4184_/S vssd1 vssd1 vccd1 vccd1 _4172_/A sky130_fd_sc_hd__mux2_1
X_3122_ _4554_/S _3158_/A _3112_/X _5287_/A _3121_/X vssd1 vssd1 vccd1 vccd1 _3122_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4248__A2 _4228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3053_ _3053_/A _3288_/C _3053_/C _3052_/A vssd1 vssd1 vccd1 vccd1 _3054_/A sky130_fd_sc_hd__or4b_1
XFILLER_67_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5599__A _6104_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_304 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3955_ _3996_/B vssd1 vssd1 vccd1 vccd1 _3983_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4956__B1 _3723_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2906_ _3824_/A _6005_/Q vssd1 vssd1 vccd1 vccd1 _3315_/B sky130_fd_sc_hd__xor2_1
XFILLER_31_370 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3886_ _3886_/A _3886_/B vssd1 vssd1 vccd1 vccd1 _3886_/Y sky130_fd_sc_hd__nor2_1
X_5625_ _5642_/B vssd1 vssd1 vccd1 vccd1 _5635_/B sky130_fd_sc_hd__clkbuf_1
X_2837_ _6008_/Q vssd1 vssd1 vccd1 vccd1 _5277_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5556_ _5597_/A vssd1 vssd1 vccd1 vccd1 _5556_/X sky130_fd_sc_hd__clkbuf_2
X_4507_ _4518_/D _4504_/Y _4506_/Y _4460_/X vssd1 vssd1 vccd1 vccd1 _5860_/D sky130_fd_sc_hd__o211a_1
X_5487_ _6063_/Q _5490_/B vssd1 vssd1 vccd1 vccd1 _5487_/X sky130_fd_sc_hd__or2_1
X_4438_ _4438_/A _4438_/B vssd1 vssd1 vccd1 vccd1 _4438_/X sky130_fd_sc_hd__or2_1
XFILLER_86_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4369_ _4369_/A vssd1 vssd1 vccd1 vccd1 _5826_/D sky130_fd_sc_hd__clkbuf_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5436__A1 _5357_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6108_ _6108_/CLK _6108_/D vssd1 vssd1 vccd1 vccd1 _6108_/Q sky130_fd_sc_hd__dfxtp_1
X_6039_ _6112_/CLK _6039_/D vssd1 vssd1 vccd1 vccd1 _6039_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3998__A1 _3938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4478__A2 _4331_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_454 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3740_ _5376_/A _5697_/Q _3753_/S vssd1 vssd1 vccd1 vccd1 _3741_/B sky130_fd_sc_hd__mux2_1
X_3671_ _3671_/A vssd1 vssd1 vccd1 vccd1 _5678_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5410_ _3587_/X _5404_/X _5407_/X _5409_/X vssd1 vssd1 vccd1 vccd1 _6033_/D sky130_fd_sc_hd__o211a_1
X_5341_ _5341_/A vssd1 vssd1 vccd1 vccd1 _6016_/D sky130_fd_sc_hd__clkbuf_1
X_5272_ _3867_/X _5304_/B _3066_/B _3373_/B vssd1 vssd1 vccd1 vccd1 _5272_/X sky130_fd_sc_hd__a211o_1
XANTENNA__4469__A2 _3061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4223_ _3335_/C _3938_/A _4222_/X vssd1 vssd1 vccd1 vccd1 _4447_/D sky130_fd_sc_hd__a21o_1
X_4154_ _5788_/Q _4152_/X _4167_/S vssd1 vssd1 vccd1 vccd1 _4155_/A sky130_fd_sc_hd__mux2_1
X_3105_ _4287_/A vssd1 vssd1 vccd1 vccd1 _4231_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4085_ _4085_/A vssd1 vssd1 vccd1 vccd1 _5768_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3036_ _3858_/A vssd1 vssd1 vccd1 vccd1 _3037_/A sky130_fd_sc_hd__buf_2
XFILLER_55_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_462 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4987_ _4986_/B _4982_/B _4972_/A _5928_/Q vssd1 vssd1 vccd1 vccd1 _4988_/C sky130_fd_sc_hd__a31o_1
X_3938_ _3938_/A _3938_/B vssd1 vssd1 vccd1 vccd1 _3954_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__3296__B _3296_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3869_ _3869_/A _3899_/A vssd1 vssd1 vccd1 vccd1 _3869_/X sky130_fd_sc_hd__or2_1
X_5608_ _3598_/X _5602_/X _5607_/X _5597_/X vssd1 vssd1 vccd1 vccd1 _6106_/D sky130_fd_sc_hd__o211a_1
XANTENNA__3904__A1 _3287_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5539_ _6081_/Q _5549_/B vssd1 vssd1 vccd1 vccd1 _5539_/X sky130_fd_sc_hd__or2_1
XFILLER_11_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_15_wb_clk_i clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6014_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_86_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4396__A1 _5834_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput17 la_data_in[43] vssd1 vssd1 vccd1 vccd1 _5389_/A sky130_fd_sc_hd__clkbuf_1
Xinput28 la_data_in[53] vssd1 vssd1 vccd1 vccd1 _3611_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_10_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput39 la_data_in[63] vssd1 vssd1 vccd1 vccd1 _5075_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_6_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3950__A _3966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4320__A1 _3275_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output51_A _5878_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4084__A0 _5768_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5890_ _5892_/CLK _5890_/D vssd1 vssd1 vccd1 vccd1 _5890_/Q sky130_fd_sc_hd__dfxtp_1
X_4910_ _4870_/X _4908_/X _4909_/X _4875_/X vssd1 vssd1 vccd1 vccd1 _4910_/X sky130_fd_sc_hd__o211a_1
X_4841_ _6112_/Q _4840_/X _4873_/S vssd1 vssd1 vccd1 vccd1 _4841_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4772_ _6081_/Q _4783_/B vssd1 vssd1 vccd1 vccd1 _4772_/X sky130_fd_sc_hd__or2_1
XFILLER_20_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3723_ _5876_/Q _5875_/Q _3723_/C _3722_/X vssd1 vssd1 vccd1 vccd1 _3724_/A sky130_fd_sc_hd__or4b_1
XANTENNA__5336__A0 _6067_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3654_ _3738_/A _5174_/A vssd1 vssd1 vccd1 vccd1 _3678_/S sky130_fd_sc_hd__nand2_1
X_3585_ _5295_/A vssd1 vssd1 vccd1 vccd1 _3585_/X sky130_fd_sc_hd__clkbuf_2
X_5324_ _5309_/A _5315_/B _5281_/B _5321_/Y vssd1 vssd1 vccd1 vccd1 _5324_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5639__A1 _5366_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5255_ _5255_/A _5255_/B vssd1 vssd1 vccd1 vccd1 _5255_/X sky130_fd_sc_hd__or2_1
X_4206_ _4206_/A _4455_/A _3379_/A vssd1 vssd1 vccd1 vccd1 _4206_/X sky130_fd_sc_hd__or3b_1
XFILLER_68_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5186_ _5186_/A _5186_/B vssd1 vssd1 vccd1 vccd1 _5187_/A sky130_fd_sc_hd__and2_1
XFILLER_28_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4167__S _4167_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4137_ _5783_/Q _4135_/X _4150_/S vssd1 vssd1 vccd1 vccd1 _4138_/A sky130_fd_sc_hd__mux2_1
X_4068_ _4068_/A vssd1 vssd1 vccd1 vccd1 _5763_/D sky130_fd_sc_hd__clkbuf_1
X_3019_ _5285_/A _3407_/A _3469_/C _3432_/B _5301_/B vssd1 vssd1 vccd1 vccd1 _3019_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3100__A _3135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3586__C1 _3585_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3889__A0 _3869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_40 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3370_ _6131_/Q vssd1 vssd1 vccd1 vccd1 _4455_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _5944_/Q _5038_/A _5039_/Y vssd1 vssd1 vccd1 vccd1 _5944_/D sky130_fd_sc_hd__o21a_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5942_ _5942_/CLK _5942_/D vssd1 vssd1 vccd1 vccd1 _5942_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3839__B _3839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3804__B1 _3525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3280__A1 _5336_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5873_ _5988_/CLK _5873_/D vssd1 vssd1 vccd1 vccd1 _5873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4016__A _4113_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4824_ _4824_/A vssd1 vssd1 vccd1 vccd1 _4824_/X sky130_fd_sc_hd__clkbuf_2
X_4755_ _5891_/Q _4705_/X _4753_/X _4754_/X vssd1 vssd1 vccd1 vccd1 _5891_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3706_ _3706_/A vssd1 vssd1 vccd1 vccd1 _5688_/D sky130_fd_sc_hd__clkbuf_1
X_4686_ _6024_/Q _4674_/X _4675_/X vssd1 vssd1 vccd1 vccd1 _4686_/X sky130_fd_sc_hd__o21a_1
X_3637_ _3637_/A vssd1 vssd1 vccd1 vccd1 _5668_/D sky130_fd_sc_hd__clkbuf_1
X_3568_ _4881_/A vssd1 vssd1 vccd1 vccd1 _5624_/A sky130_fd_sc_hd__buf_2
X_5307_ _5307_/A _5307_/B _5294_/S vssd1 vssd1 vccd1 vccd1 _5307_/X sky130_fd_sc_hd__or3b_1
XFILLER_88_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3499_ _3357_/X _3505_/C _3496_/Y _3498_/X _4322_/A vssd1 vssd1 vccd1 vccd1 _6123_/D
+ sky130_fd_sc_hd__a32o_1
X_5238_ _5238_/A vssd1 vssd1 vccd1 vccd1 _6005_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5169_ _5391_/A vssd1 vssd1 vccd1 vccd1 _5169_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_29_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4048__A0 _6100_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_40_wb_clk_i_A clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__4599__A1 _4717_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3765__A _3765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3484__B _3484_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_30_wb_clk_i clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5942_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4596__A _6065_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2870_ _5814_/Q vssd1 vssd1 vccd1 vccd1 _3044_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_15_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4540_ _4541_/A _4541_/B vssd1 vssd1 vccd1 vccd1 _4542_/B sky130_fd_sc_hd__nor2_1
Xuser_proj_example_273 vssd1 vssd1 vccd1 vccd1 io_out[21] user_proj_example_273/LO
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_262 vssd1 vssd1 vccd1 vccd1 io_out[10] user_proj_example_262/LO
+ sky130_fd_sc_hd__conb_1
X_4471_ _4471_/A _4471_/B vssd1 vssd1 vccd1 vccd1 _4471_/Y sky130_fd_sc_hd__nor2_1
Xuser_proj_example_251 vssd1 vssd1 vccd1 vccd1 user_proj_example_251/HI wbs_dat_o[30]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_240 vssd1 vssd1 vccd1 vccd1 user_proj_example_240/HI wbs_dat_o[19]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_284 vssd1 vssd1 vccd1 vccd1 io_out[32] user_proj_example_284/LO
+ sky130_fd_sc_hd__conb_1
X_3422_ _3076_/Y _3266_/Y _3085_/X _3117_/B vssd1 vssd1 vccd1 vccd1 _3423_/D sky130_fd_sc_hd__o211a_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ _3161_/A _3335_/X _3352_/X _4458_/A vssd1 vssd1 vccd1 vccd1 _3353_/X sky130_fd_sc_hd__o211a_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3284_ _3117_/B _3886_/A _4470_/B vssd1 vssd1 vccd1 vccd1 _3284_/Y sky130_fd_sc_hd__o21ai_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6072_ _6118_/CLK _6072_/D vssd1 vssd1 vccd1 vccd1 _6072_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5023_ _5939_/Q _5938_/Q _5023_/C vssd1 vssd1 vccd1 vccd1 _5030_/C sky130_fd_sc_hd__and3_1
XFILLER_65_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5925_ _5988_/CLK _5925_/D vssd1 vssd1 vccd1 vccd1 _5925_/Q sky130_fd_sc_hd__dfxtp_1
X_5856_ _6014_/CLK _5856_/D vssd1 vssd1 vccd1 vccd1 _5856_/Q sky130_fd_sc_hd__dfxtp_1
X_4807_ _4858_/A vssd1 vssd1 vccd1 vccd1 _4807_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2999_ _5719_/Q _4471_/A vssd1 vssd1 vccd1 vccd1 _3891_/A sky130_fd_sc_hd__nor2_1
XANTENNA__4180__S _4184_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5787_ _6048_/CLK _5787_/D vssd1 vssd1 vccd1 vccd1 _5787_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3585__A _5295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4753__A1 _6055_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4738_ _6138_/Q _4737_/X _4770_/S vssd1 vssd1 vccd1 vccd1 _4738_/X sky130_fd_sc_hd__mux2_1
X_4669_ _6071_/Q _4683_/B vssd1 vssd1 vccd1 vccd1 _4669_/X sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_7_wb_clk_i_A _5813_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5466__C1 _5461_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3492__B2 _3491_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3492__A1 _3505_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_368 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4680__A0 _6120_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3971_ _3971_/A vssd1 vssd1 vccd1 vccd1 _5728_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4432__A0 _5975_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2922_ _2949_/C vssd1 vssd1 vccd1 vccd1 _2959_/C sky130_fd_sc_hd__clkbuf_2
X_5710_ _6087_/CLK _5710_/D vssd1 vssd1 vccd1 vccd1 _5710_/Q sky130_fd_sc_hd__dfxtp_1
X_2853_ _3272_/B _3518_/A _2853_/C _4234_/B vssd1 vssd1 vccd1 vccd1 _3127_/A sky130_fd_sc_hd__or4_1
X_5641_ _5369_/X _5623_/A _5640_/X _5638_/X vssd1 vssd1 vccd1 vccd1 _6119_/D sky130_fd_sc_hd__o211a_1
XANTENNA__4735__A1 _6029_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5572_ _5363_/X _5559_/X _5570_/X _5571_/X vssd1 vssd1 vccd1 vccd1 _6093_/D sky130_fd_sc_hd__o211a_1
X_4523_ _3146_/B _5864_/Q _4523_/S vssd1 vssd1 vccd1 vccd1 _4524_/B sky130_fd_sc_hd__mux2_1
X_4454_ _4454_/A vssd1 vssd1 vccd1 vccd1 _5848_/D sky130_fd_sc_hd__clkbuf_1
X_3405_ _3405_/A _3899_/A vssd1 vssd1 vccd1 vccd1 _3405_/X sky130_fd_sc_hd__or2_1
X_4385_ _5831_/Q _4384_/X _4391_/S vssd1 vssd1 vccd1 vccd1 _4386_/A sky130_fd_sc_hd__mux2_1
X_6124_ _6130_/CLK _6124_/D vssd1 vssd1 vccd1 vccd1 _6124_/Q sky130_fd_sc_hd__dfxtp_1
X_3336_ _5856_/Q _3481_/B vssd1 vssd1 vccd1 vccd1 _3336_/X sky130_fd_sc_hd__or2_1
XFILLER_58_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6055_ _6080_/CLK _6055_/D vssd1 vssd1 vccd1 vccd1 _6055_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3267_ _3839_/A _3928_/A vssd1 vssd1 vccd1 vccd1 _3800_/A sky130_fd_sc_hd__nor2_1
X_5006_ _5934_/Q _5933_/Q _5006_/C vssd1 vssd1 vccd1 vccd1 _5008_/A sky130_fd_sc_hd__and3_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3474__B2 _3287_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3198_ _5942_/Q vssd1 vssd1 vccd1 vccd1 _3198_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5908_ _6087_/CLK _5908_/D vssd1 vssd1 vccd1 vccd1 _5908_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5839_ _6112_/CLK _5839_/D vssd1 vssd1 vccd1 vccd1 _5839_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4726__A1 _5888_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input13_A la_data_in[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4114__A _4182_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4170_ _4170_/A vssd1 vssd1 vccd1 vccd1 _4184_/S sky130_fd_sc_hd__buf_2
X_3121_ _3161_/A _3938_/A _3117_/Y _3118_/Y _3374_/A vssd1 vssd1 vccd1 vccd1 _3121_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_67_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3052_ _3052_/A vssd1 vssd1 vccd1 vccd1 _3841_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_82_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_187 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3954_ _3954_/A _3954_/B vssd1 vssd1 vccd1 vccd1 _3996_/B sky130_fd_sc_hd__nor2_1
X_2905_ _4280_/A vssd1 vssd1 vccd1 vccd1 _3824_/A sky130_fd_sc_hd__clkbuf_4
X_3885_ _4466_/A _3901_/A vssd1 vssd1 vccd1 vccd1 _3886_/B sky130_fd_sc_hd__nand2_1
X_2836_ _5256_/B vssd1 vssd1 vccd1 vccd1 _3508_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5624_ _5624_/A _5624_/B vssd1 vssd1 vccd1 vccd1 _5642_/B sky130_fd_sc_hd__nor2_1
XANTENNA__5381__A1 _5376_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5555_ _6088_/Q _5555_/B vssd1 vssd1 vccd1 vccd1 _5555_/X sky130_fd_sc_hd__or2_1
X_4506_ _4518_/D _4506_/B vssd1 vssd1 vccd1 vccd1 _4506_/Y sky130_fd_sc_hd__nand2_1
X_5486_ _3611_/X _5470_/A _5485_/X _5477_/X vssd1 vssd1 vccd1 vccd1 _6062_/D sky130_fd_sc_hd__o211a_1
X_4437_ _4470_/A _4437_/B vssd1 vssd1 vccd1 vccd1 _4437_/Y sky130_fd_sc_hd__nor2_1
XFILLER_86_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input5_A la_data_in[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4368_ _5826_/Q _4367_/X _4374_/S vssd1 vssd1 vccd1 vccd1 _4369_/A sky130_fd_sc_hd__mux2_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4892__A0 _5959_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6107_ _6108_/CLK _6107_/D vssd1 vssd1 vccd1 vccd1 _6107_/Q sky130_fd_sc_hd__dfxtp_1
X_3319_ _3316_/X _3318_/X _3046_/A vssd1 vssd1 vccd1 vccd1 _3319_/X sky130_fd_sc_hd__a21o_1
X_4299_ _5810_/Q _4313_/C vssd1 vssd1 vccd1 vccd1 _4300_/B sky130_fd_sc_hd__xnor2_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3447__B2 _3880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3447__A1 _3857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6038_ _6112_/CLK _6038_/D vssd1 vssd1 vccd1 vccd1 _6038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3013__A _3841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4938__A1 _6040_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3670_ _3684_/A _3670_/B vssd1 vssd1 vccd1 vccd1 _3671_/A sky130_fd_sc_hd__and2_1
XFILLER_40_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5340_ _6016_/Q _5339_/X _5340_/S vssd1 vssd1 vccd1 vccd1 _5341_/A sky130_fd_sc_hd__mux2_1
X_5271_ _5277_/B _5271_/B vssd1 vssd1 vccd1 vccd1 _5271_/Y sky130_fd_sc_hd__xnor2_1
X_4222_ _6124_/Q _5714_/Q _5836_/Q _6129_/Q vssd1 vssd1 vccd1 vccd1 _4222_/X sky130_fd_sc_hd__a22o_1
X_4153_ _4170_/A vssd1 vssd1 vccd1 vccd1 _4167_/S sky130_fd_sc_hd__buf_2
XFILLER_83_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3104_ _5250_/A vssd1 vssd1 vccd1 vccd1 _4287_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4084_ _5768_/Q _4082_/X _4097_/S vssd1 vssd1 vccd1 vccd1 _4085_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3035_ _3858_/A _3837_/A _3035_/C vssd1 vssd1 vccd1 vccd1 _3035_/X sky130_fd_sc_hd__and3_1
XFILLER_63_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4986_ _5928_/Q _4986_/B _5855_/Q _5016_/D vssd1 vssd1 vccd1 vccd1 _4993_/C sky130_fd_sc_hd__and4_1
X_3937_ _4236_/A _3936_/X _5847_/Q vssd1 vssd1 vccd1 vccd1 _3938_/B sky130_fd_sc_hd__o21a_1
XFILLER_11_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3868_ _3869_/A _3079_/B _3849_/C _5761_/Q vssd1 vssd1 vccd1 vccd1 _3868_/X sky130_fd_sc_hd__a31o_1
XFILLER_31_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3799_ _3799_/A vssd1 vssd1 vccd1 vccd1 _5713_/D sky130_fd_sc_hd__clkbuf_1
X_5607_ _6106_/Q _5614_/B vssd1 vssd1 vccd1 vccd1 _5607_/X sky130_fd_sc_hd__or2_1
XFILLER_11_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5538_ _5555_/B vssd1 vssd1 vccd1 vccd1 _5549_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_87_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5469_ _5601_/A _5469_/B vssd1 vssd1 vccd1 vccd1 _5470_/A sky130_fd_sc_hd__or2_1
XFILLER_74_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_55_wb_clk_i clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _5703_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_14_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5042__B1 _3135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5593__A1 _5393_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput18 la_data_in[44] vssd1 vssd1 vccd1 vccd1 _5393_/A sky130_fd_sc_hd__clkbuf_1
Xinput29 la_data_in[54] vssd1 vssd1 vccd1 vccd1 _3614_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__5223__A _5295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4840_ _5665_/Q _4839_/X _4872_/S vssd1 vssd1 vccd1 vccd1 _4840_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4771_ _6105_/Q _4770_/X _4771_/S vssd1 vssd1 vccd1 vccd1 _4771_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5584__A1 _5376_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3722_ input8/X _5692_/Q _3722_/S vssd1 vssd1 vccd1 vccd1 _3722_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3653_ _3653_/A vssd1 vssd1 vccd1 vccd1 _5673_/D sky130_fd_sc_hd__clkbuf_1
X_5323_ _5323_/A _5323_/B vssd1 vssd1 vccd1 vccd1 _5323_/X sky130_fd_sc_hd__or2_1
X_3584_ _5544_/A vssd1 vssd1 vccd1 vccd1 _5295_/A sky130_fd_sc_hd__clkbuf_4
X_5254_ _5254_/A _5254_/B _5254_/C _5254_/D vssd1 vssd1 vccd1 vccd1 _5260_/B sky130_fd_sc_hd__or4_1
X_4205_ _4205_/A vssd1 vssd1 vccd1 vccd1 _5248_/B sky130_fd_sc_hd__inv_2
XANTENNA__3860__B _3897_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5185_ _5062_/A _5992_/Q _5189_/S vssd1 vssd1 vccd1 vccd1 _5186_/B sky130_fd_sc_hd__mux2_1
X_4136_ _4170_/A vssd1 vssd1 vccd1 vccd1 _4150_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_83_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_30_wb_clk_i_A clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4067_ _5763_/Q _4065_/X _4080_/S vssd1 vssd1 vccd1 vccd1 _4068_/A sky130_fd_sc_hd__mux2_1
X_3018_ _3297_/B vssd1 vssd1 vccd1 vccd1 _3432_/B sky130_fd_sc_hd__clkinv_2
XANTENNA__3822__B2 _3331_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4969_ _4982_/C _4975_/B _4955_/X vssd1 vssd1 vccd1 vccd1 _4970_/C sky130_fd_sc_hd__o21ai_1
XFILLER_22_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5941_ _5941_/CLK _5941_/D vssd1 vssd1 vccd1 vccd1 _5941_/Q sky130_fd_sc_hd__dfxtp_1
X_5872_ _6131_/CLK _5872_/D vssd1 vssd1 vccd1 vccd1 _5872_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3280__A2 _3255_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_0_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6135_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_4823_ _6086_/Q _4834_/B vssd1 vssd1 vccd1 vccd1 _4823_/X sky130_fd_sc_hd__or2_1
XFILLER_33_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4754_ _6031_/Q _4744_/X _4745_/X vssd1 vssd1 vccd1 vccd1 _4754_/X sky130_fd_sc_hd__o21a_1
X_3705_ _3732_/A _3705_/B vssd1 vssd1 vccd1 vccd1 _3706_/A sky130_fd_sc_hd__and2_1
X_4685_ _6048_/Q _4654_/X _4664_/X _4684_/X vssd1 vssd1 vccd1 vccd1 _4685_/X sky130_fd_sc_hd__a211o_1
XANTENNA__4032__A _4203_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3636_ _3648_/A _3636_/B vssd1 vssd1 vccd1 vccd1 _3637_/A sky130_fd_sc_hd__and2_1
X_3567_ _3712_/B _4604_/A vssd1 vssd1 vccd1 vccd1 _4881_/A sky130_fd_sc_hd__or2_1
XFILLER_88_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5306_ _5302_/X _5305_/X _4041_/S vssd1 vssd1 vccd1 vccd1 _5307_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_458 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3498_ _3354_/X _3522_/B _3497_/X _3412_/X vssd1 vssd1 vccd1 vccd1 _3498_/X sky130_fd_sc_hd__a31o_1
X_5237_ _5232_/X _3480_/B _5237_/S vssd1 vssd1 vccd1 vccd1 _5238_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5168_ _5986_/Q _5168_/B vssd1 vssd1 vccd1 vccd1 _5168_/X sky130_fd_sc_hd__or2_1
XFILLER_56_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3810__S _5278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4906__S _4914_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5099_ _5072_/X _5080_/A _5097_/X _5098_/X vssd1 vssd1 vccd1 vccd1 _5961_/D sky130_fd_sc_hd__o211a_1
X_4119_ _4170_/A vssd1 vssd1 vccd1 vccd1 _4133_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_16_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5548__A1 _3604_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3731__A0 _5369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input43_A wbs_sel_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4596__B _4917_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xuser_proj_example_230 vssd1 vssd1 vccd1 vccd1 user_proj_example_230/HI wbs_dat_o[9]
+ sky130_fd_sc_hd__conb_1
XFILLER_30_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_proj_example_263 vssd1 vssd1 vccd1 vccd1 io_out[11] user_proj_example_263/LO
+ sky130_fd_sc_hd__conb_1
X_4470_ _4470_/A _4470_/B _4470_/C vssd1 vssd1 vccd1 vccd1 _4470_/X sky130_fd_sc_hd__and3_1
Xuser_proj_example_252 vssd1 vssd1 vccd1 vccd1 user_proj_example_252/HI wbs_dat_o[31]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_241 vssd1 vssd1 vccd1 vccd1 user_proj_example_241/HI wbs_dat_o[20]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_285 vssd1 vssd1 vccd1 vccd1 io_out[33] user_proj_example_285/LO
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_274 vssd1 vssd1 vccd1 vccd1 io_out[22] user_proj_example_274/LO
+ sky130_fd_sc_hd__conb_1
X_3421_ _3522_/A vssd1 vssd1 vccd1 vccd1 _3505_/C sky130_fd_sc_hd__clkbuf_2
X_3352_ _3508_/B _3928_/B _3348_/X _3351_/X vssd1 vssd1 vccd1 vccd1 _3352_/X sky130_fd_sc_hd__a211o_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3722__A0 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3283_ _3838_/A _3283_/B vssd1 vssd1 vccd1 vccd1 _4470_/B sky130_fd_sc_hd__nor2_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6071_ _6118_/CLK _6071_/D vssd1 vssd1 vccd1 vccd1 _6071_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5022_ _5938_/Q _5023_/C _5021_/Y vssd1 vssd1 vccd1 vccd1 _5938_/D sky130_fd_sc_hd__a21oi_1
XFILLER_78_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5411__A _6034_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5924_ _5988_/CLK _5924_/D vssd1 vssd1 vccd1 vccd1 _5924_/Q sky130_fd_sc_hd__dfxtp_1
X_5855_ _5945_/CLK _5855_/D vssd1 vssd1 vccd1 vccd1 _5855_/Q sky130_fd_sc_hd__dfxtp_1
X_4806_ _5896_/Q _4756_/X _4802_/X _4805_/X vssd1 vssd1 vccd1 vccd1 _5896_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2998_ _3481_/B vssd1 vssd1 vccd1 vccd1 _4471_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5786_ _6048_/CLK _5786_/D vssd1 vssd1 vccd1 vccd1 _5786_/Q sky130_fd_sc_hd__dfxtp_1
X_4737_ _5702_/Q _5679_/Q _4748_/S vssd1 vssd1 vccd1 vccd1 _4737_/X sky130_fd_sc_hd__mux2_1
X_4668_ _6095_/Q _4667_/X _4668_/S vssd1 vssd1 vccd1 vccd1 _4668_/X sky130_fd_sc_hd__mux2_1
X_3619_ _3617_/X _3592_/A _3618_/X _3609_/X vssd1 vssd1 vccd1 vccd1 _5665_/D sky130_fd_sc_hd__o211a_1
X_4599_ _4717_/A _4593_/X _4596_/X _5469_/B vssd1 vssd1 vccd1 vccd1 _4599_/X sky130_fd_sc_hd__o211a_1
XFILLER_88_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2945__A _4218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4636__S _4645_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_406 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3970_ _3994_/A _3970_/B vssd1 vssd1 vccd1 vccd1 _3971_/A sky130_fd_sc_hd__and2_1
XFILLER_62_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2921_ _2933_/A vssd1 vssd1 vccd1 vccd1 _3429_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3686__A _4251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2852_ _3118_/B _2852_/B vssd1 vssd1 vccd1 vccd1 _4234_/B sky130_fd_sc_hd__nand2_1
X_5640_ _6119_/Q _5642_/B vssd1 vssd1 vccd1 vccd1 _5640_/X sky130_fd_sc_hd__or2_1
X_5571_ _5597_/A vssd1 vssd1 vccd1 vccd1 _5571_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4522_ _5857_/Q _4568_/B _3542_/A _4480_/Y vssd1 vssd1 vccd1 vccd1 _4523_/S sky130_fd_sc_hd__a22o_1
X_4453_ _4524_/A _4453_/B vssd1 vssd1 vccd1 vccd1 _4454_/A sky130_fd_sc_hd__and2_1
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3404_ _3842_/A _3800_/A vssd1 vssd1 vccd1 vccd1 _3899_/A sky130_fd_sc_hd__nand2_1
X_4384_ _6053_/Q _5830_/Q _4396_/S vssd1 vssd1 vccd1 vccd1 _4384_/X sky130_fd_sc_hd__mux2_1
X_3335_ _5256_/A _5258_/A _3335_/C _4236_/A vssd1 vssd1 vccd1 vccd1 _3335_/X sky130_fd_sc_hd__or4_1
X_6123_ _6130_/CLK _6123_/D vssd1 vssd1 vccd1 vccd1 _6123_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3266_ _3266_/A _3898_/A vssd1 vssd1 vccd1 vccd1 _3266_/Y sky130_fd_sc_hd__nor2_1
X_6054_ _6080_/CLK _6054_/D vssd1 vssd1 vccd1 vccd1 _6054_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5005_ _5005_/A _5005_/B vssd1 vssd1 vccd1 vccd1 _5933_/D sky130_fd_sc_hd__nor2_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3474__A2 _3869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3197_ _5016_/D vssd1 vssd1 vccd1 vccd1 _4954_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_53_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5907_ _6003_/CLK _5907_/D vssd1 vssd1 vccd1 vccd1 _5907_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4191__S _4200_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5838_ _5941_/CLK _5838_/D vssd1 vssd1 vccd1 vccd1 _5838_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5769_ _5914_/CLK _5769_/D vssd1 vssd1 vccd1 vccd1 _5769_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4220__A _4220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4874__B _4885_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4662__A1 _6022_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6032__D _6032_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5226__A _5295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3120_ _5243_/B vssd1 vssd1 vccd1 vccd1 _3374_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_67_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3051_ _5851_/Q vssd1 vssd1 vccd1 vccd1 _3052_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_67_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4405__A1 _6060_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3953_ _3953_/A vssd1 vssd1 vccd1 vccd1 _3953_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2904_ _5848_/Q vssd1 vssd1 vccd1 vccd1 _4280_/A sky130_fd_sc_hd__clkbuf_2
X_3884_ _6104_/Q _3882_/X _4041_/S vssd1 vssd1 vccd1 vccd1 _3884_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2835_ _3335_/C vssd1 vssd1 vccd1 vccd1 _5256_/B sky130_fd_sc_hd__clkbuf_1
X_5623_ _5623_/A vssd1 vssd1 vccd1 vccd1 _5623_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5554_ _3614_/X _5536_/A _5553_/X _5545_/X vssd1 vssd1 vccd1 vccd1 _6087_/D sky130_fd_sc_hd__o211a_1
X_4505_ _4511_/A vssd1 vssd1 vccd1 vccd1 _4506_/B sky130_fd_sc_hd__inv_2
X_5485_ _6062_/Q _5490_/B vssd1 vssd1 vccd1 vccd1 _5485_/X sky130_fd_sc_hd__or2_1
X_4436_ _4436_/A _4450_/D vssd1 vssd1 vccd1 vccd1 _4436_/Y sky130_fd_sc_hd__nor2_1
X_4367_ _6048_/Q _5825_/Q _4380_/S vssd1 vssd1 vccd1 vccd1 _4367_/X sky130_fd_sc_hd__mux2_1
X_3318_ _4437_/B _3432_/B _2983_/B _3469_/C _3046_/B vssd1 vssd1 vccd1 vccd1 _3318_/X
+ sky130_fd_sc_hd__o2111a_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6106_ _6108_/CLK _6106_/D vssd1 vssd1 vccd1 vccd1 _6106_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4298_ _4315_/A _4313_/C _4298_/C vssd1 vssd1 vccd1 vccd1 _5809_/D sky130_fd_sc_hd__nor3_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2926__C _4438_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3249_ _4436_/A vssd1 vssd1 vccd1 vccd1 _5171_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_73_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6037_ _6064_/CLK _6037_/D vssd1 vssd1 vccd1 vccd1 _6037_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4644__A1 _5880_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4914__S _4914_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3907__B1 _5775_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4096__S _4110_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4635__A1 _5879_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3013__B _3839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4399__A0 _6059_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5270_ _3373_/B _3066_/B _5278_/D _5269_/X vssd1 vssd1 vccd1 vccd1 _5274_/A sky130_fd_sc_hd__o22a_1
XANTENNA__3126__B2 _3547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4221_ _5256_/A _3081_/B _3355_/X vssd1 vssd1 vccd1 vccd1 _4447_/C sky130_fd_sc_hd__a21o_1
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4152_ _6138_/Q _5787_/Q _4162_/S vssd1 vssd1 vccd1 vccd1 _4152_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3103_ _4218_/A vssd1 vssd1 vccd1 vccd1 _5250_/A sky130_fd_sc_hd__clkbuf_2
X_4083_ _4203_/S vssd1 vssd1 vccd1 vccd1 _4097_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__5403__B _5403_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_20_wb_clk_i_A _5836_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3034_ _5721_/Q vssd1 vssd1 vccd1 vccd1 _3858_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_55_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3204__A _6022_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4985_ _4985_/A vssd1 vssd1 vccd1 vccd1 _5927_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3936_ _5240_/A _5287_/B _3936_/C vssd1 vssd1 vccd1 vccd1 _3936_/X sky130_fd_sc_hd__or3_1
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3867_ _3867_/A vssd1 vssd1 vccd1 vccd1 _3867_/X sky130_fd_sc_hd__clkbuf_2
X_3798_ input5/X _5343_/B _3798_/C _4607_/A vssd1 vssd1 vccd1 vccd1 _3799_/A sky130_fd_sc_hd__and4_1
X_5606_ _3587_/X _5602_/X _5605_/X _5597_/X vssd1 vssd1 vccd1 vccd1 _6105_/D sky130_fd_sc_hd__o211a_1
X_5537_ _5603_/A _5537_/B vssd1 vssd1 vccd1 vccd1 _5555_/B sky130_fd_sc_hd__nor2_1
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5468_ _3582_/X _5449_/A _5467_/X _5461_/X vssd1 vssd1 vccd1 vccd1 _6056_/D sky130_fd_sc_hd__o211a_1
X_5399_ _6031_/Q _5399_/B vssd1 vssd1 vccd1 vccd1 _5399_/X sky130_fd_sc_hd__or2_1
X_4419_ _5971_/Q _5841_/Q _4426_/S vssd1 vssd1 vccd1 vccd1 _4419_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_24_wb_clk_i clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5988_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_3_3__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput19 la_data_in[45] vssd1 vssd1 vccd1 vccd1 _5396_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_10_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4856__A1 _5979_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4608__A1 _6017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4554__S _4554_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5569__C1 _5556_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4770_ _5658_/Q _4769_/X _4770_/S vssd1 vssd1 vccd1 vccd1 _4770_/X sky130_fd_sc_hd__mux2_1
X_3721_ _4575_/A _3720_/X _3999_/A vssd1 vssd1 vccd1 vccd1 _5691_/D sky130_fd_sc_hd__a21oi_1
XFILLER_9_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3652_ _3666_/A _3652_/B vssd1 vssd1 vccd1 vccd1 _3653_/A sky130_fd_sc_hd__and2_1
X_3583_ _5657_/Q _5648_/B vssd1 vssd1 vccd1 vccd1 _3583_/X sky130_fd_sc_hd__or2_1
X_5322_ _5315_/A _5315_/B _5321_/Y vssd1 vssd1 vccd1 vccd1 _5322_/X sky130_fd_sc_hd__a21o_1
XFILLER_5_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5253_ _4241_/A _5278_/B _4555_/C _4288_/A _3832_/A vssd1 vssd1 vccd1 vccd1 _5254_/D
+ sky130_fd_sc_hd__a2111o_1
X_4204_ _4204_/A vssd1 vssd1 vccd1 vccd1 _5803_/D sky130_fd_sc_hd__clkbuf_1
X_5184_ _5184_/A vssd1 vssd1 vccd1 vccd1 _5991_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4135_ _6133_/Q _3037_/A _4145_/S vssd1 vssd1 vccd1 vccd1 _4135_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5272__A1 _3867_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3869__A _3869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4066_ _4203_/S vssd1 vssd1 vccd1 vccd1 _4080_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_83_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3017_ _3853_/C _3017_/B vssd1 vssd1 vccd1 vccd1 _3469_/C sky130_fd_sc_hd__or2_1
XFILLER_43_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4968_ _5923_/Q _4968_/B _4968_/C vssd1 vssd1 vccd1 vccd1 _4975_/B sky130_fd_sc_hd__and3_1
XFILLER_11_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3586__A1 _3582_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3919_ _5782_/Q _3916_/X _3918_/X _3460_/C _2858_/A vssd1 vssd1 vccd1 vccd1 _3919_/X
+ sky130_fd_sc_hd__a221o_1
X_4899_ _5952_/Q _4898_/X _4915_/S vssd1 vssd1 vccd1 vccd1 _4899_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3109__A _5234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5234__A _5234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5940_ _5942_/CLK _5940_/D vssd1 vssd1 vccd1 vccd1 _5940_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3804__A2 _3379_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5871_ _6005_/CLK _5871_/D vssd1 vssd1 vccd1 vccd1 _5871_/Q sky130_fd_sc_hd__dfxtp_1
X_4822_ _6110_/Q _4821_/X _4822_/S vssd1 vssd1 vccd1 vccd1 _4822_/X sky130_fd_sc_hd__mux2_1
X_4753_ _6055_/Q _4706_/X _4716_/X _4752_/X vssd1 vssd1 vccd1 vccd1 _4753_/X sky130_fd_sc_hd__a211o_1
XFILLER_21_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3704_ _3614_/A _5688_/Q _3707_/S vssd1 vssd1 vccd1 vccd1 _3705_/B sky130_fd_sc_hd__mux2_1
XANTENNA__5409__A _5461_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4684_ _4665_/X _4682_/X _4683_/X _4670_/X vssd1 vssd1 vccd1 vccd1 _4684_/X sky130_fd_sc_hd__o211a_1
X_3635_ input7/X _5668_/Q _3641_/S vssd1 vssd1 vccd1 vccd1 _3636_/B sky130_fd_sc_hd__mux2_1
X_3566_ _3711_/A _4594_/B vssd1 vssd1 vccd1 vccd1 _4604_/A sky130_fd_sc_hd__or2_1
X_5305_ _5246_/B _5299_/Y _5303_/X _5304_/Y _3867_/X vssd1 vssd1 vccd1 vccd1 _5305_/X
+ sky130_fd_sc_hd__o221a_1
X_3497_ _5255_/A vssd1 vssd1 vccd1 vccd1 _3497_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5236_ _5261_/A _5236_/B _5236_/C _5236_/D vssd1 vssd1 vccd1 vccd1 _5237_/S sky130_fd_sc_hd__or4_1
XFILLER_56_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5167_ _5072_/X _5149_/A _5166_/X _5158_/X vssd1 vssd1 vccd1 vccd1 _5985_/D sky130_fd_sc_hd__o211a_1
XFILLER_68_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5098_ _5141_/A vssd1 vssd1 vccd1 vccd1 _5098_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4118_ _6115_/Q _5777_/Q _4128_/S vssd1 vssd1 vccd1 vccd1 _4118_/X sky130_fd_sc_hd__mux2_1
X_4049_ _4203_/S vssd1 vssd1 vccd1 vccd1 _4063_/S sky130_fd_sc_hd__buf_2
XANTENNA__4577__D_N _3564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4194__S _4200_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3822__A1_N _3071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input36_A la_data_in[60] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_proj_example_220 vssd1 vssd1 vccd1 vccd1 user_proj_example_220/HI la_data_out[127]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_264 vssd1 vssd1 vccd1 vccd1 io_out[12] user_proj_example_264/LO
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_253 vssd1 vssd1 vccd1 vccd1 io_oeb[1] user_proj_example_253/LO
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_242 vssd1 vssd1 vccd1 vccd1 user_proj_example_242/HI wbs_dat_o[21]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_231 vssd1 vssd1 vccd1 vccd1 user_proj_example_231/HI wbs_dat_o[10]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_286 vssd1 vssd1 vccd1 vccd1 io_out[34] user_proj_example_286/LO
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_275 vssd1 vssd1 vccd1 vccd1 io_out[23] user_proj_example_275/LO
+ sky130_fd_sc_hd__conb_1
X_3420_ _5171_/A _3420_/B vssd1 vssd1 vccd1 vccd1 _5855_/D sky130_fd_sc_hd__nor2_1
X_3351_ _3349_/X _3520_/A _3410_/A vssd1 vssd1 vccd1 vccd1 _3351_/X sky130_fd_sc_hd__o21a_1
XANTENNA__3722__A1 _5692_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3282_ _3282_/A _3282_/B vssd1 vssd1 vccd1 vccd1 _3886_/A sky130_fd_sc_hd__nand2_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6070_ _6091_/CLK _6070_/D vssd1 vssd1 vccd1 vccd1 _6070_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5021_ _5938_/Q _5023_/C _5020_/X vssd1 vssd1 vccd1 vccd1 _5021_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_26_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3212__A _6021_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5923_ _5988_/CLK _5923_/D vssd1 vssd1 vccd1 vccd1 _5923_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5854_ _5988_/CLK _5854_/D vssd1 vssd1 vccd1 vccd1 _5854_/Q sky130_fd_sc_hd__dfxtp_1
X_4805_ _6036_/Q _4803_/X _4804_/X vssd1 vssd1 vccd1 vccd1 _4805_/X sky130_fd_sc_hd__o21a_1
X_2997_ _2997_/A vssd1 vssd1 vccd1 vccd1 _3481_/B sky130_fd_sc_hd__clkbuf_2
X_5785_ _6138_/CLK _5785_/D vssd1 vssd1 vccd1 vccd1 _5785_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4736_ _5889_/Q _4705_/X _4734_/X _4735_/X vssd1 vssd1 vccd1 vccd1 _5889_/D sky130_fd_sc_hd__a22o_1
X_4667_ _6119_/Q _4666_/X _4667_/S vssd1 vssd1 vccd1 vccd1 _4667_/X sky130_fd_sc_hd__mux2_1
X_3618_ _5665_/Q _3618_/B vssd1 vssd1 vccd1 vccd1 _3618_/X sky130_fd_sc_hd__or2_1
X_4598_ _5126_/A vssd1 vssd1 vccd1 vccd1 _5469_/B sky130_fd_sc_hd__buf_2
X_3549_ _3546_/Y _3547_/Y _3548_/X _5740_/Q _3255_/X vssd1 vssd1 vccd1 vccd1 _5740_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5466__A1 _3563_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5219_ _5069_/A _6002_/Q _5225_/S vssd1 vssd1 vccd1 vccd1 _5220_/B sky130_fd_sc_hd__mux2_1
XFILLER_84_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5049__A _5622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3792__A _3966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4099__S _4110_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5457__A1 _5386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_418 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3032__A _3897_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2920_ _6009_/Q _6008_/Q _6007_/Q _6006_/Q vssd1 vssd1 vccd1 vccd1 _2933_/A sky130_fd_sc_hd__nand4b_1
XFILLER_62_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2851_ _3049_/A _5736_/Q vssd1 vssd1 vccd1 vccd1 _2852_/B sky130_fd_sc_hd__nand2_1
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5570_ _6093_/Q _5570_/B vssd1 vssd1 vccd1 vccd1 _5570_/X sky130_fd_sc_hd__or2_1
X_4521_ _4521_/A vssd1 vssd1 vccd1 vccd1 _5863_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4452_ _3354_/X _4449_/X _4452_/S vssd1 vssd1 vccd1 vccd1 _4453_/B sky130_fd_sc_hd__mux2_1
X_3403_ _5715_/Q vssd1 vssd1 vccd1 vccd1 _3405_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4383_ _4383_/A vssd1 vssd1 vccd1 vccd1 _4396_/S sky130_fd_sc_hd__clkbuf_4
X_6122_ _6122_/CLK _6122_/D vssd1 vssd1 vccd1 vccd1 _6122_/Q sky130_fd_sc_hd__dfxtp_1
X_3334_ _6123_/Q _6126_/Q _6130_/Q _6129_/Q vssd1 vssd1 vccd1 vccd1 _4236_/A sky130_fd_sc_hd__or4_2
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3265_ _3854_/A vssd1 vssd1 vccd1 vccd1 _3898_/A sky130_fd_sc_hd__clkbuf_2
X_6053_ _6080_/CLK _6053_/D vssd1 vssd1 vccd1 vccd1 _6053_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5422__A _6039_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5004_ _5933_/Q _5006_/C _4990_/X vssd1 vssd1 vccd1 vccd1 _5005_/B sky130_fd_sc_hd__o21ai_1
XFILLER_38_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3196_ _3196_/A _3196_/B _3196_/C vssd1 vssd1 vccd1 vccd1 _5016_/D sky130_fd_sc_hd__nor3_1
XFILLER_81_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3631__A0 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5906_ _5986_/CLK _5906_/D vssd1 vssd1 vccd1 vccd1 _5906_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5837_ _5941_/CLK _5837_/D vssd1 vssd1 vccd1 vccd1 _5837_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5768_ _5941_/CLK _5768_/D vssd1 vssd1 vccd1 vccd1 _5768_/Q sky130_fd_sc_hd__dfxtp_1
X_4719_ _6136_/Q _4718_/X _4719_/S vssd1 vssd1 vccd1 vccd1 _4719_/X sky130_fd_sc_hd__mux2_1
X_5699_ _6080_/CLK _5699_/D vssd1 vssd1 vccd1 vccd1 _5699_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_49_wb_clk_i clkbuf_3_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6088_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_89_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3787__A _5188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3050_ _3853_/A vssd1 vssd1 vccd1 vccd1 _5241_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4405__A2 _3802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3952_ _3952_/A vssd1 vssd1 vccd1 vccd1 _3953_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2903_ _3873_/D vssd1 vssd1 vccd1 vccd1 _4255_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3883_ _4231_/A vssd1 vssd1 vccd1 vccd1 _4041_/S sky130_fd_sc_hd__clkbuf_4
X_2834_ _6128_/Q vssd1 vssd1 vccd1 vccd1 _3335_/C sky130_fd_sc_hd__clkbuf_2
X_5622_ _5622_/A _5622_/B vssd1 vssd1 vccd1 vccd1 _5623_/A sky130_fd_sc_hd__or2_1
XANTENNA__3377__C1 _3525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5553_ _6087_/Q _5555_/B vssd1 vssd1 vccd1 vccd1 _5553_/X sky130_fd_sc_hd__or2_1
X_4504_ _4511_/A _4504_/B vssd1 vssd1 vccd1 vccd1 _4504_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5417__A _6037_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5484_ _3607_/X _5470_/X _5483_/X _5477_/X vssd1 vssd1 vccd1 vccd1 _6061_/D sky130_fd_sc_hd__o211a_1
X_4435_ _3936_/X _4003_/X _4001_/Y vssd1 vssd1 vccd1 vccd1 _4450_/D sky130_fd_sc_hd__o21ai_1
XFILLER_6_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4366_ _4366_/A vssd1 vssd1 vccd1 vccd1 _4380_/S sky130_fd_sc_hd__clkbuf_2
X_3317_ _3317_/A vssd1 vssd1 vccd1 vccd1 _4437_/B sky130_fd_sc_hd__clkbuf_2
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6105_ _6108_/CLK _6105_/D vssd1 vssd1 vccd1 vccd1 _6105_/Q sky130_fd_sc_hd__dfxtp_1
X_4297_ _5809_/Q _4297_/B vssd1 vssd1 vccd1 vccd1 _4298_/C sky130_fd_sc_hd__nor2_1
XANTENNA__5152__A _5979_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3248_ _5011_/A vssd1 vssd1 vccd1 vccd1 _4436_/A sky130_fd_sc_hd__buf_2
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6036_ _6088_/CLK _6036_/D vssd1 vssd1 vccd1 vccd1 _6036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3179_ _5924_/Q _4939_/A _5913_/Q _3174_/Y _3178_/X vssd1 vssd1 vccd1 vccd1 _3196_/A
+ sky130_fd_sc_hd__a221o_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3907__A1 _5255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4885__B _4885_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5062__A _5062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4571__B2 _5875_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4220_ _4220_/A _4220_/B vssd1 vssd1 vccd1 vccd1 _4220_/Y sky130_fd_sc_hd__nor2_1
X_4151_ _4151_/A vssd1 vssd1 vccd1 vccd1 _5787_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3102_ _4002_/A vssd1 vssd1 vccd1 vccd1 _4218_/A sky130_fd_sc_hd__clkbuf_2
X_4082_ _6111_/Q _5767_/Q _4092_/S vssd1 vssd1 vccd1 vccd1 _4082_/X sky130_fd_sc_hd__mux2_1
X_3033_ _3031_/Y _3032_/X _5301_/A vssd1 vssd1 vccd1 vccd1 _3059_/B sky130_fd_sc_hd__o21bai_1
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4984_ _4995_/B _4984_/B _4984_/C vssd1 vssd1 vccd1 vccd1 _4985_/A sky130_fd_sc_hd__and3_1
X_3935_ _4218_/A _6124_/Q _3935_/C _6121_/Q vssd1 vssd1 vccd1 vccd1 _3936_/C sky130_fd_sc_hd__or4_1
XFILLER_51_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5339__A0 _6068_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3866_ _3866_/A vssd1 vssd1 vccd1 vccd1 _5717_/D sky130_fd_sc_hd__clkbuf_1
X_5605_ _6105_/Q _5614_/B vssd1 vssd1 vccd1 vccd1 _5605_/X sky130_fd_sc_hd__or2_1
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3797_ _4855_/A vssd1 vssd1 vccd1 vccd1 _4607_/A sky130_fd_sc_hd__clkbuf_2
X_5536_ _5536_/A vssd1 vssd1 vccd1 vccd1 _5536_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5467_ _6056_/Q _5467_/B vssd1 vssd1 vccd1 vccd1 _5467_/X sky130_fd_sc_hd__or2_1
X_4418_ _4418_/A vssd1 vssd1 vccd1 vccd1 _5841_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5398_ _5396_/X _5387_/B _5397_/X _5391_/X vssd1 vssd1 vccd1 vccd1 _6030_/D sky130_fd_sc_hd__o211a_1
X_4349_ _4366_/A vssd1 vssd1 vccd1 vccd1 _4363_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__4197__S _4200_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5275__C1 _5169_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6019_ _6067_/CLK _6019_/D vssd1 vssd1 vccd1 vccd1 _6019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4553__A1 _3454_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4305__A1 _3275_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4136__A _4170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3720_ _5875_/Q _3719_/X vssd1 vssd1 vccd1 vccd1 _3720_/X sky130_fd_sc_hd__or2b_1
XFILLER_9_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3651_ _5373_/A _5673_/Q _3651_/S vssd1 vssd1 vccd1 vccd1 _3652_/B sky130_fd_sc_hd__mux2_1
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3582_ _3582_/A vssd1 vssd1 vccd1 vccd1 _3582_/X sky130_fd_sc_hd__buf_2
X_5321_ _5327_/A vssd1 vssd1 vccd1 vccd1 _5321_/Y sky130_fd_sc_hd__inv_2
X_5252_ _5252_/A _5252_/B vssd1 vssd1 vccd1 vccd1 _5278_/B sky130_fd_sc_hd__nor2_2
X_4203_ _5803_/Q _4202_/X _4203_/S vssd1 vssd1 vccd1 vccd1 _4204_/A sky130_fd_sc_hd__mux2_1
X_5183_ _5186_/A _5183_/B vssd1 vssd1 vccd1 vccd1 _5184_/A sky130_fd_sc_hd__and2_1
X_4134_ _4134_/A vssd1 vssd1 vccd1 vccd1 _5782_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4065_ _6106_/Q _5762_/Q _4075_/S vssd1 vssd1 vccd1 vccd1 _4065_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5430__A _6041_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3016_ _4255_/A _2863_/A _3428_/B _3430_/A _5301_/A vssd1 vssd1 vccd1 vccd1 _3016_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4967_ _4968_/B _4948_/A _4968_/C _5923_/Q vssd1 vssd1 vccd1 vccd1 _4970_/B sky130_fd_sc_hd__a31o_1
XANTENNA__3885__A _4466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3918_ _3037_/A _3917_/Y _4322_/B _3463_/X _5782_/Q vssd1 vssd1 vccd1 vccd1 _3918_/X
+ sky130_fd_sc_hd__a32o_1
X_4898_ _6002_/Q _5994_/Q _4898_/S vssd1 vssd1 vccd1 vccd1 _4898_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3849_ _3849_/A _3849_/B _3849_/C vssd1 vssd1 vccd1 vccd1 _3901_/B sky130_fd_sc_hd__and3_1
X_5519_ _5376_/X _5514_/X _5517_/X _5518_/X vssd1 vssd1 vccd1 vccd1 _6073_/D sky130_fd_sc_hd__o211a_1
XANTENNA__5605__A _6105_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_44 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2964__A _3038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4390__S _4396_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3723__D_N _3722_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5515__A _5581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5250__A _5250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5870_ _5874_/CLK _5870_/D vssd1 vssd1 vccd1 vccd1 _5870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4821_ _5663_/Q _4820_/X _4821_/S vssd1 vssd1 vccd1 vccd1 _4821_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4214__B1 _3296_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4752_ _4717_/X _4750_/X _4751_/X _4722_/X vssd1 vssd1 vccd1 vccd1 _4752_/X sky130_fd_sc_hd__o211a_1
XANTENNA__4765__A1 _5401_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3703_ _3770_/A vssd1 vssd1 vccd1 vccd1 _3732_/A sky130_fd_sc_hd__clkbuf_2
X_4683_ _6072_/Q _4683_/B vssd1 vssd1 vccd1 vccd1 _4683_/X sky130_fd_sc_hd__or2_1
X_3634_ _3668_/A vssd1 vssd1 vccd1 vccd1 _3648_/A sky130_fd_sc_hd__clkbuf_1
X_3565_ input3/X input2/X input4/X vssd1 vssd1 vccd1 vccd1 _4594_/B sky130_fd_sc_hd__or3_2
XFILLER_88_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5304_ _5304_/A _5304_/B vssd1 vssd1 vccd1 vccd1 _5304_/Y sky130_fd_sc_hd__nor2_1
X_3496_ _3496_/A _3496_/B vssd1 vssd1 vccd1 vccd1 _3496_/Y sky130_fd_sc_hd__nor2_1
XFILLER_88_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5235_ _3901_/A _5234_/Y _4555_/B _5254_/A vssd1 vssd1 vccd1 vccd1 _5236_/D sky130_fd_sc_hd__a211o_1
X_5166_ _5985_/Q _5168_/B vssd1 vssd1 vccd1 vccd1 _5166_/X sky130_fd_sc_hd__or2_1
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4117_ _4117_/A vssd1 vssd1 vccd1 vccd1 _5777_/D sky130_fd_sc_hd__clkbuf_1
X_5097_ _5961_/Q _5100_/B vssd1 vssd1 vccd1 vccd1 _5097_/X sky130_fd_sc_hd__or2_1
X_4048_ _6100_/Q _5757_/Q _4058_/S vssd1 vssd1 vccd1 vccd1 _4048_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3008__A1 _3842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5999_ _5999_/CLK _5999_/D vssd1 vssd1 vccd1 vccd1 _5999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4893__B _4917_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input29_A la_data_in[54] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_316 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4747__A1 _5890_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_proj_example_210 vssd1 vssd1 vccd1 vccd1 user_proj_example_210/HI la_data_out[117]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_221 vssd1 vssd1 vccd1 vccd1 user_proj_example_221/HI wbs_dat_o[0]
+ sky130_fd_sc_hd__conb_1
XFILLER_11_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xuser_proj_example_254 vssd1 vssd1 vccd1 vccd1 io_out[2] user_proj_example_254/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_7_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuser_proj_example_243 vssd1 vssd1 vccd1 vccd1 user_proj_example_243/HI wbs_dat_o[22]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_232 vssd1 vssd1 vccd1 vccd1 user_proj_example_232/HI wbs_dat_o[11]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_287 vssd1 vssd1 vccd1 vccd1 io_out[35] user_proj_example_287/LO
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_276 vssd1 vssd1 vccd1 vccd1 io_out[24] user_proj_example_276/LO
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_265 vssd1 vssd1 vccd1 vccd1 io_out[13] user_proj_example_265/LO
+ sky130_fd_sc_hd__conb_1
X_3350_ _3350_/A _3350_/B _3350_/C vssd1 vssd1 vccd1 vccd1 _3520_/A sky130_fd_sc_hd__and3_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ _5025_/B vssd1 vssd1 vccd1 vccd1 _5020_/X sky130_fd_sc_hd__clkbuf_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3281_ _5717_/Q vssd1 vssd1 vccd1 vccd1 _3282_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5922_ _5922_/CLK _5922_/D vssd1 vssd1 vccd1 vccd1 _5922_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5853_ _5945_/CLK _5853_/D vssd1 vssd1 vccd1 vccd1 _5853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5784_ _6138_/CLK _5784_/D vssd1 vssd1 vccd1 vccd1 _5784_/Q sky130_fd_sc_hd__dfxtp_1
X_4804_ _4855_/A vssd1 vssd1 vccd1 vccd1 _4804_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2996_ _5848_/Q _5719_/Q vssd1 vssd1 vccd1 vccd1 _3297_/B sky130_fd_sc_hd__xor2_1
X_4735_ _6029_/Q _4674_/X _4675_/X vssd1 vssd1 vccd1 vccd1 _4735_/X sky130_fd_sc_hd__o21a_1
X_4666_ _5695_/Q _5672_/Q _4697_/S vssd1 vssd1 vccd1 vccd1 _4666_/X sky130_fd_sc_hd__mux2_1
X_4597_ _4597_/A _4604_/B vssd1 vssd1 vccd1 vccd1 _5126_/A sky130_fd_sc_hd__or2_1
X_3617_ _3617_/A vssd1 vssd1 vccd1 vccd1 _3617_/X sky130_fd_sc_hd__clkbuf_2
X_3548_ _4548_/A _5859_/Q _3540_/X _3544_/C _5858_/Q vssd1 vssd1 vccd1 vccd1 _3548_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_88_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3479_ _3046_/A _3470_/X _3472_/X _3478_/X vssd1 vssd1 vccd1 vccd1 _3479_/X sky130_fd_sc_hd__o211a_1
X_5218_ _5218_/A vssd1 vssd1 vccd1 vccd1 _6001_/D sky130_fd_sc_hd__clkbuf_1
X_5149_ _5149_/A vssd1 vssd1 vccd1 vccd1 _5149_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4426__A0 _5973_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4218__B _4218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3229__B2 _5387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3313__A _3326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2850_ _3038_/A vssd1 vssd1 vccd1 vccd1 _3049_/A sky130_fd_sc_hd__buf_2
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4520_ _4524_/A _4520_/B vssd1 vssd1 vccd1 vccd1 _4521_/A sky130_fd_sc_hd__and2_1
X_4451_ _5847_/Q _4436_/Y _4449_/X _4450_/X vssd1 vssd1 vccd1 vccd1 _5847_/D sky130_fd_sc_hd__o22a_1
X_3402_ _5715_/Q vssd1 vssd1 vccd1 vccd1 _3402_/Y sky130_fd_sc_hd__inv_2
X_6121_ _6121_/CLK _6121_/D vssd1 vssd1 vccd1 vccd1 _6121_/Q sky130_fd_sc_hd__dfxtp_1
X_4382_ _4382_/A vssd1 vssd1 vccd1 vccd1 _5830_/D sky130_fd_sc_hd__clkbuf_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3333_ _6124_/Q vssd1 vssd1 vccd1 vccd1 _5258_/A sky130_fd_sc_hd__clkbuf_2
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3264_ _3264_/A vssd1 vssd1 vccd1 vccd1 _3854_/A sky130_fd_sc_hd__clkbuf_2
X_6052_ _6080_/CLK _6052_/D vssd1 vssd1 vccd1 vccd1 _6052_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5003_ _5933_/Q _5006_/C vssd1 vssd1 vccd1 vccd1 _5005_/A sky130_fd_sc_hd__and2_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3195_ _4953_/A _5910_/Q _3186_/Y _3188_/X _3194_/X vssd1 vssd1 vccd1 vccd1 _3196_/C
+ sky130_fd_sc_hd__a2111o_1
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3631__A1 _5667_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5905_ _5999_/CLK _5905_/D vssd1 vssd1 vccd1 vccd1 _5905_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5836_ _5836_/CLK _5836_/D vssd1 vssd1 vccd1 vccd1 _5836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2979_ _2975_/Y _4217_/A _4220_/A _3440_/A vssd1 vssd1 vccd1 vccd1 _3300_/A sky130_fd_sc_hd__and4bb_1
X_5767_ _5941_/CLK _5767_/D vssd1 vssd1 vccd1 vccd1 _5767_/Q sky130_fd_sc_hd__dfxtp_1
X_4718_ _5700_/Q _5677_/Q _4748_/S vssd1 vssd1 vccd1 vccd1 _4718_/X sky130_fd_sc_hd__mux2_1
X_5698_ _6080_/CLK _5698_/D vssd1 vssd1 vccd1 vccd1 _5698_/Q sky130_fd_sc_hd__dfxtp_1
X_4649_ _4611_/X _4647_/X _4648_/X _4620_/X vssd1 vssd1 vccd1 vccd1 _4649_/X sky130_fd_sc_hd__o211a_1
XANTENNA__3117__B _3117_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_18_wb_clk_i _5836_/CLK vssd1 vssd1 vccd1 vccd1 _6130_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_84_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2972__A _3256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5375__A1 _5373_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_6_wb_clk_i_A clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_90_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3951_ _3951_/A vssd1 vssd1 vccd1 vccd1 _5724_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2902_ _5814_/Q _5817_/Q _2949_/D _5815_/Q vssd1 vssd1 vccd1 vccd1 _3873_/D sky130_fd_sc_hd__or4bb_2
XFILLER_50_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3613__A1 _3611_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3882_ _3867_/X _3868_/X _3869_/X _3881_/X _5761_/Q vssd1 vssd1 vccd1 vccd1 _3882_/X
+ sky130_fd_sc_hd__a32o_1
X_2833_ _3053_/C vssd1 vssd1 vccd1 vccd1 _3518_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5621_ _3617_/X _5602_/A _5620_/X _5612_/X vssd1 vssd1 vccd1 vccd1 _6112_/D sky130_fd_sc_hd__o211a_1
X_5552_ _3611_/X _5536_/A _5551_/X _5545_/X vssd1 vssd1 vccd1 vccd1 _6086_/D sky130_fd_sc_hd__o211a_1
XANTENNA__4602__A _4716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4503_ _4529_/A _3146_/B _4562_/A vssd1 vssd1 vccd1 vccd1 _4504_/B sky130_fd_sc_hd__a21oi_1
X_5483_ _6061_/Q _5483_/B vssd1 vssd1 vccd1 vccd1 _5483_/X sky130_fd_sc_hd__or2_1
X_4434_ _4434_/A vssd1 vssd1 vccd1 vccd1 _5846_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4365_ _4365_/A vssd1 vssd1 vccd1 vccd1 _5825_/D sky130_fd_sc_hd__clkbuf_1
X_3316_ _3428_/A _3314_/X _3315_/Y _3448_/A vssd1 vssd1 vccd1 vccd1 _3316_/X sky130_fd_sc_hd__a211o_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6104_ _6135_/CLK _6104_/D vssd1 vssd1 vccd1 vccd1 _6104_/Q sky130_fd_sc_hd__dfxtp_1
X_4296_ _5809_/Q _4297_/B vssd1 vssd1 vccd1 vccd1 _4313_/C sky130_fd_sc_hd__and2_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6035_ _6108_/CLK _6035_/D vssd1 vssd1 vccd1 vccd1 _6035_/Q sky130_fd_sc_hd__dfxtp_1
X_3247_ _5873_/Q vssd1 vssd1 vccd1 vccd1 _3247_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4049__A _4203_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3178_ _4968_/B _4935_/A _4931_/A _5920_/Q vssd1 vssd1 vccd1 vccd1 _3178_/X sky130_fd_sc_hd__a22o_1
XFILLER_26_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5819_ _6117_/CLK _5819_/D vssd1 vssd1 vccd1 vccd1 _5819_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4512__A _5284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5327__B _5327_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4317__C1 _3867_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input11_A la_data_in[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3798__A input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4393__S _4396_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5518__A _5529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3038__A _3038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4150_ _5787_/Q _4149_/X _4150_/S vssd1 vssd1 vccd1 vccd1 _4151_/A sky130_fd_sc_hd__mux2_1
X_3101_ _6122_/Q vssd1 vssd1 vccd1 vccd1 _4002_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_68_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4081_ _4081_/A vssd1 vssd1 vccd1 vccd1 _5767_/D sky130_fd_sc_hd__clkbuf_1
X_3032_ _3897_/A _4283_/A _3494_/B _3304_/B vssd1 vssd1 vccd1 vccd1 _3032_/X sky130_fd_sc_hd__and4_1
XFILLER_55_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4983_ _4982_/B _4982_/C _4986_/B vssd1 vssd1 vccd1 vccd1 _4984_/C sky130_fd_sc_hd__a21o_1
XFILLER_51_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5587__A1 _5382_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3934_ _5252_/A vssd1 vssd1 vccd1 vccd1 _5287_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3865_ _3282_/A _3823_/X _3865_/S vssd1 vssd1 vccd1 vccd1 _3866_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4332__A _4399_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5428__A _5471_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5604_ _5620_/B vssd1 vssd1 vccd1 vccd1 _5614_/B sky130_fd_sc_hd__clkbuf_1
X_3796_ input3/X _4577_/B input2/X _3564_/B vssd1 vssd1 vccd1 vccd1 _4855_/A sky130_fd_sc_hd__nor4b_4
X_5535_ _5601_/A _5535_/B vssd1 vssd1 vccd1 vccd1 _5536_/A sky130_fd_sc_hd__or2_1
X_5466_ _3563_/X _5449_/A _5465_/X _5461_/X vssd1 vssd1 vccd1 vccd1 _6055_/D sky130_fd_sc_hd__o211a_1
X_4417_ _5841_/Q _4416_/X _4417_/S vssd1 vssd1 vccd1 vccd1 _4418_/A sky130_fd_sc_hd__mux2_1
X_5397_ _6030_/Q _5399_/B vssd1 vssd1 vccd1 vccd1 _5397_/X sky130_fd_sc_hd__or2_1
XFILLER_86_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input3_A la_data_in[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4348_ _4348_/A vssd1 vssd1 vccd1 vccd1 _5820_/D sky130_fd_sc_hd__clkbuf_1
X_4279_ _3423_/A _3081_/B _4278_/X vssd1 vssd1 vccd1 vccd1 _4279_/X sky130_fd_sc_hd__o21ba_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6018_ _6018_/CLK _6018_/D vssd1 vssd1 vccd1 vccd1 _6018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5578__A1 _5373_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4553__A2 _3326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4305__A2 _3497_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_33_wb_clk_i clkbuf_3_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6112_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_77_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5569__A1 _5360_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3650_ _3668_/A vssd1 vssd1 vccd1 vccd1 _3666_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3581_ _3563_/X _3576_/X _3580_/X _3221_/X vssd1 vssd1 vccd1 vccd1 _5656_/D sky130_fd_sc_hd__o211a_1
X_5320_ _5320_/A _5320_/B vssd1 vssd1 vccd1 vccd1 _5320_/Y sky130_fd_sc_hd__nand2_1
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5251_ _5287_/A _5251_/B _5278_/C _5268_/B vssd1 vssd1 vccd1 vccd1 _5251_/X sky130_fd_sc_hd__or4b_1
XFILLER_5_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4202_ _5953_/Q _5802_/Q _4554_/S vssd1 vssd1 vccd1 vccd1 _4202_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5182_ _5059_/A _5991_/Q _5189_/S vssd1 vssd1 vccd1 vccd1 _5183_/B sky130_fd_sc_hd__mux2_1
X_4133_ _5782_/Q _4132_/X _4133_/S vssd1 vssd1 vccd1 vccd1 _4134_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4064_ _4064_/A vssd1 vssd1 vccd1 vccd1 _5762_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3015_ _3015_/A vssd1 vssd1 vccd1 vccd1 _5301_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4327__A _4327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3231__A _6033_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4966_ _4966_/A _4966_/B _4966_/C vssd1 vssd1 vccd1 vccd1 _5922_/D sky130_fd_sc_hd__nor3_1
X_3917_ _3917_/A vssd1 vssd1 vccd1 vccd1 _3917_/Y sky130_fd_sc_hd__inv_2
X_4897_ _5905_/Q _4858_/X _4895_/X _4896_/X vssd1 vssd1 vccd1 vccd1 _5905_/D sky130_fd_sc_hd__a22o_1
XANTENNA__5158__A _5391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3848_ _5254_/A _4555_/B _4555_/C _5261_/A vssd1 vssd1 vccd1 vccd1 _3913_/A sky130_fd_sc_hd__or4_1
X_3779_ _3779_/A vssd1 vssd1 vccd1 vccd1 _5708_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5518_ _5529_/A vssd1 vssd1 vccd1 vccd1 _5518_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5449_ _5449_/A vssd1 vssd1 vccd1 vccd1 _5449_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_23 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3141__A _3408_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4038__B1_N _3821_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5515__B _5535_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3986__A _3999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2890__A _3159_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4820_ _5710_/Q _5687_/Q _4848_/S vssd1 vssd1 vccd1 vccd1 _4820_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3422__C1 _3117_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4751_ _6079_/Q _4783_/B vssd1 vssd1 vccd1 vccd1 _4751_/X sky130_fd_sc_hd__or2_1
X_3702_ _3702_/A vssd1 vssd1 vccd1 vccd1 _5687_/D sky130_fd_sc_hd__clkbuf_1
X_4682_ _6096_/Q _4680_/X _4720_/S vssd1 vssd1 vccd1 vccd1 _4682_/X sky130_fd_sc_hd__mux2_1
X_3633_ _3633_/A vssd1 vssd1 vccd1 vccd1 _5667_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3725__A0 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3564_ _4580_/A _3564_/B vssd1 vssd1 vccd1 vccd1 _3712_/B sky130_fd_sc_hd__nand2_1
XANTENNA__4610__A _4716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5303_ _5297_/A _5243_/B _3424_/B _5304_/B vssd1 vssd1 vccd1 vccd1 _5303_/X sky130_fd_sc_hd__o211a_1
X_3495_ _3493_/X _3274_/C _4239_/B _3494_/Y _3396_/Y vssd1 vssd1 vccd1 vccd1 _3496_/B
+ sky130_fd_sc_hd__o221a_1
X_5234_ _5234_/A _5234_/B vssd1 vssd1 vccd1 vccd1 _5234_/Y sky130_fd_sc_hd__nor2_1
X_5165_ _5069_/X _5149_/A _5164_/X _5158_/X vssd1 vssd1 vccd1 vccd1 _5984_/D sky130_fd_sc_hd__o211a_1
XFILLER_68_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4116_ _5777_/Q _4115_/X _4116_/S vssd1 vssd1 vccd1 vccd1 _4117_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5096_ _5069_/X _5080_/A _5095_/X _5087_/X vssd1 vssd1 vccd1 vccd1 _5960_/D sky130_fd_sc_hd__o211a_1
XFILLER_83_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4047_ _4047_/A vssd1 vssd1 vccd1 vccd1 _5757_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5998_ _5999_/CLK _5998_/D vssd1 vssd1 vccd1 vccd1 _5998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4949_ _5855_/Q _5854_/Q _5853_/Q vssd1 vssd1 vccd1 vccd1 _4964_/B sky130_fd_sc_hd__or3_1
XFILLER_24_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3716__A0 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3136__A _3547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2975__A _3826_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5351__A _6017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_proj_example_211 vssd1 vssd1 vccd1 vccd1 user_proj_example_211/HI la_data_out[118]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_200 vssd1 vssd1 vccd1 vccd1 user_proj_example_200/HI la_data_out[107]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_255 vssd1 vssd1 vccd1 vccd1 io_out[3] user_proj_example_255/LO
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_233 vssd1 vssd1 vccd1 vccd1 user_proj_example_233/HI wbs_dat_o[12]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_244 vssd1 vssd1 vccd1 vccd1 user_proj_example_244/HI wbs_dat_o[23]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_222 vssd1 vssd1 vccd1 vccd1 user_proj_example_222/HI wbs_dat_o[1]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_288 vssd1 vssd1 vccd1 vccd1 io_out[36] user_proj_example_288/LO
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_277 vssd1 vssd1 vccd1 vccd1 io_out[25] user_proj_example_277/LO
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_266 vssd1 vssd1 vccd1 vccd1 io_out[14] user_proj_example_266/LO
+ sky130_fd_sc_hd__conb_1
X_3280_ _5336_/S _3255_/X _3271_/X _3272_/Y _3279_/X vssd1 vssd1 vccd1 vccd1 _6132_/D
+ sky130_fd_sc_hd__a32o_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4132__A0 _6119_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2885__A _3071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5921_ _5922_/CLK _5921_/D vssd1 vssd1 vccd1 vccd1 _5921_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5852_ _5988_/CLK _5852_/D vssd1 vssd1 vccd1 vccd1 _5852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5783_ _6048_/CLK _5783_/D vssd1 vssd1 vccd1 vccd1 _5783_/Q sky130_fd_sc_hd__dfxtp_1
X_4803_ _5403_/B vssd1 vssd1 vccd1 vccd1 _4803_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2995_ _3845_/C vssd1 vssd1 vccd1 vccd1 _3440_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4734_ _6053_/Q _4706_/X _4716_/X _4733_/X vssd1 vssd1 vccd1 vccd1 _4734_/X sky130_fd_sc_hd__a211o_1
X_4665_ _4717_/A vssd1 vssd1 vccd1 vccd1 _4665_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4596_ _6065_/Q _4917_/B vssd1 vssd1 vccd1 vccd1 _4596_/X sky130_fd_sc_hd__or2_1
X_3616_ _3614_/X _3592_/A _3615_/X _3609_/X vssd1 vssd1 vccd1 vccd1 _5664_/D sky130_fd_sc_hd__o211a_1
X_3547_ _3547_/A _3556_/A vssd1 vssd1 vccd1 vccd1 _3547_/Y sky130_fd_sc_hd__nor2_1
X_3478_ _3475_/X _3477_/X _3484_/A vssd1 vssd1 vccd1 vccd1 _3478_/X sky130_fd_sc_hd__a21o_1
XFILLER_69_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5217_ _5220_/A _5217_/B vssd1 vssd1 vccd1 vccd1 _5218_/A sky130_fd_sc_hd__and2_1
XANTENNA__5171__A _5171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5148_ _5405_/B _5148_/B vssd1 vssd1 vccd1 vccd1 _5149_/A sky130_fd_sc_hd__or2_1
XFILLER_28_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5079_ _5601_/B _5148_/B vssd1 vssd1 vccd1 vccd1 _5080_/A sky130_fd_sc_hd__or2_1
XFILLER_71_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4515__A _4970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4250__A _4276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3165__B2 _3071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input41_A wbs_cyc_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4396__S _4396_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5081__A _5603_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3032__C _3494_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4450_ _5011_/A _4450_/B _5287_/B _4450_/D vssd1 vssd1 vccd1 vccd1 _4450_/X sky130_fd_sc_hd__or4_1
X_3401_ _3423_/B _3802_/B _3502_/A vssd1 vssd1 vccd1 vccd1 _3496_/A sky130_fd_sc_hd__or3_1
X_4381_ _5830_/Q _4380_/X _4391_/S vssd1 vssd1 vccd1 vccd1 _4382_/A sky130_fd_sc_hd__mux2_1
X_3332_ _3043_/X _3301_/X _3329_/Y _3331_/X vssd1 vssd1 vccd1 vccd1 _3332_/X sky130_fd_sc_hd__o31a_1
X_6120_ _6135_/CLK _6120_/D vssd1 vssd1 vccd1 vccd1 _6120_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3263_ _3085_/X _3509_/A _3423_/C vssd1 vssd1 vccd1 vccd1 _3263_/X sky130_fd_sc_hd__and3b_1
XFILLER_58_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6051_ _6101_/CLK _6051_/D vssd1 vssd1 vccd1 vccd1 _6051_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3194_ _3189_/Y _3190_/X _3191_/Y _3192_/X _3193_/X vssd1 vssd1 vccd1 vccd1 _3194_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ _5006_/C _5002_/B vssd1 vssd1 vccd1 vccd1 _5932_/D sky130_fd_sc_hd__nor2_1
XFILLER_26_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5904_ _5999_/CLK _5904_/D vssd1 vssd1 vccd1 vccd1 _5904_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5835_ _6014_/CLK _5835_/D vssd1 vssd1 vccd1 vccd1 _5835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2978_ _3873_/A vssd1 vssd1 vccd1 vccd1 _4220_/A sky130_fd_sc_hd__clkbuf_2
X_5766_ _6109_/CLK _5766_/D vssd1 vssd1 vccd1 vccd1 _5766_/Q sky130_fd_sc_hd__dfxtp_1
X_5697_ _6080_/CLK _5697_/D vssd1 vssd1 vccd1 vccd1 _5697_/Q sky130_fd_sc_hd__dfxtp_1
X_4717_ _4717_/A vssd1 vssd1 vccd1 vccd1 _4717_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4648_ _6069_/Q _4683_/B vssd1 vssd1 vccd1 vccd1 _4648_/X sky130_fd_sc_hd__or2_1
XANTENNA__4895__A1 _5975_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4579_ _4756_/A vssd1 vssd1 vccd1 vccd1 _4579_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_58_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6080_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_55_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5076__A _5954_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5532__C1 _5529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3950_ _3966_/A _3950_/B vssd1 vssd1 vccd1 vccd1 _3951_/A sky130_fd_sc_hd__and2_1
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2901_ _5816_/Q vssd1 vssd1 vccd1 vccd1 _2949_/D sky130_fd_sc_hd__clkbuf_1
X_3881_ _5301_/C _3880_/X _3111_/X vssd1 vssd1 vccd1 vccd1 _3881_/X sky130_fd_sc_hd__a21o_1
XFILLER_43_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2832_ _5813_/Q _2880_/A vssd1 vssd1 vccd1 vccd1 _3053_/C sky130_fd_sc_hd__or2_1
X_5620_ _6112_/Q _5620_/B vssd1 vssd1 vccd1 vccd1 _5620_/X sky130_fd_sc_hd__or2_1
X_5551_ _6086_/Q _5555_/B vssd1 vssd1 vccd1 vccd1 _5551_/X sky130_fd_sc_hd__or2_1
X_4502_ _4502_/A _4502_/B _4502_/C vssd1 vssd1 vccd1 vccd1 _4511_/A sky130_fd_sc_hd__or3_2
XFILLER_6_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5482_ _3604_/X _5470_/X _5481_/X _5477_/X vssd1 vssd1 vccd1 vccd1 _6060_/D sky130_fd_sc_hd__o211a_1
X_4433_ _5846_/Q _4432_/X _4433_/S vssd1 vssd1 vccd1 vccd1 _4434_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4877__A1 _5973_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4364_ _5825_/Q _4363_/X _4374_/S vssd1 vssd1 vccd1 vccd1 _4365_/A sky130_fd_sc_hd__mux2_1
X_3315_ _3428_/A _3315_/B vssd1 vssd1 vccd1 vccd1 _3315_/Y sky130_fd_sc_hd__nor2_1
X_4295_ _4233_/X _4297_/B _4294_/X _3723_/C vssd1 vssd1 vccd1 vccd1 _4315_/A sky130_fd_sc_hd__a31o_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6103_ _6118_/CLK _6103_/D vssd1 vssd1 vccd1 vccd1 _6103_/Q sky130_fd_sc_hd__dfxtp_1
X_3246_ _3224_/Y _4981_/B _3245_/X vssd1 vssd1 vccd1 vccd1 _5853_/D sky130_fd_sc_hd__o21a_1
XFILLER_58_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6034_ _6108_/CLK _6034_/D vssd1 vssd1 vccd1 vccd1 _6034_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3234__A _6031_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3301__A1 _4458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3177_ _5911_/Q vssd1 vssd1 vccd1 vccd1 _4931_/A sky130_fd_sc_hd__inv_2
XFILLER_81_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5818_ _6014_/CLK _5818_/D vssd1 vssd1 vccd1 vccd1 _5818_/Q sky130_fd_sc_hd__dfxtp_2
X_5749_ _5796_/CLK _5749_/D vssd1 vssd1 vccd1 vccd1 _5749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5624__A _5624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5343__B _5343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3144__A _5874_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3798__B _5343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4253__C1 _4438_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3100_ _3135_/A _3508_/C vssd1 vssd1 vccd1 vccd1 _3100_/Y sky130_fd_sc_hd__nand2_1
Xoutput80 _5907_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[94] sky130_fd_sc_hd__buf_2
X_4080_ _5767_/Q _4079_/X _4080_/S vssd1 vssd1 vccd1 vccd1 _4081_/A sky130_fd_sc_hd__mux2_1
X_3031_ _3897_/A _4283_/A _3037_/B vssd1 vssd1 vccd1 vccd1 _3031_/Y sky130_fd_sc_hd__nor3_1
XFILLER_48_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4982_ _4986_/B _4982_/B _4982_/C vssd1 vssd1 vccd1 vccd1 _4984_/B sky130_fd_sc_hd__nand3_1
XFILLER_23_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3933_ _6131_/Q _6125_/Q vssd1 vssd1 vccd1 vccd1 _5252_/A sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_3_wb_clk_i _5813_/CLK vssd1 vssd1 vccd1 vccd1 _6115_/CLK sky130_fd_sc_hd__clkbuf_16
X_3864_ _5233_/B _3888_/A vssd1 vssd1 vccd1 vccd1 _3865_/S sky130_fd_sc_hd__nor2_1
XFILLER_31_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5603_ _5603_/A _5603_/B vssd1 vssd1 vccd1 vccd1 _5620_/B sky130_fd_sc_hd__nor2_1
X_3795_ input4/X _3711_/A _4580_/A _3411_/B _5171_/B vssd1 vssd1 vccd1 vccd1 _4577_/B
+ sky130_fd_sc_hd__a311o_1
X_5534_ _3582_/X _5514_/A _5533_/X _5529_/X vssd1 vssd1 vccd1 vccd1 _6080_/D sky130_fd_sc_hd__o211a_1
X_5465_ _6055_/Q _5467_/B vssd1 vssd1 vccd1 vccd1 _5465_/X sky130_fd_sc_hd__or2_1
X_4416_ _6064_/Q _5840_/Q _4426_/S vssd1 vssd1 vccd1 vccd1 _4416_/X sky130_fd_sc_hd__mux2_1
X_5396_ _5396_/A vssd1 vssd1 vccd1 vccd1 _5396_/X sky130_fd_sc_hd__buf_2
XFILLER_59_537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4347_ _5820_/Q _4346_/X _4357_/S vssd1 vssd1 vccd1 vccd1 _4348_/A sky130_fd_sc_hd__mux2_1
X_4278_ _3335_/C _4277_/Y _3402_/Y _4235_/C vssd1 vssd1 vccd1 vccd1 _4278_/X sky130_fd_sc_hd__a22o_1
X_6017_ _6067_/CLK _6017_/D vssd1 vssd1 vccd1 vccd1 _6017_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3229_ _6032_/Q _3226_/Y _5928_/Q _5387_/A _3228_/Y vssd1 vssd1 vccd1 vccd1 _3243_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_36_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_283 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3411__B _3411_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4553__A3 _4322_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2978__A _3873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5354__A _5354_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4710__A0 _6099_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5529__A _5529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3049__A _3049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3580_ _5656_/Q _5648_/B vssd1 vssd1 vccd1 vccd1 _3580_/X sky130_fd_sc_hd__or2_1
X_5250_ _5250_/A _5256_/B _5287_/B _3502_/A vssd1 vssd1 vccd1 vccd1 _5268_/B sky130_fd_sc_hd__or4b_1
XFILLER_5_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4201_ _4201_/A vssd1 vssd1 vccd1 vccd1 _5802_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5181_ _5181_/A vssd1 vssd1 vccd1 vccd1 _5990_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4132_ _6119_/Q _5781_/Q _4145_/S vssd1 vssd1 vccd1 vccd1 _4132_/X sky130_fd_sc_hd__mux2_1
X_4063_ _5762_/Q _4062_/X _4063_/S vssd1 vssd1 vccd1 vccd1 _4064_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3014_ _3038_/A _5871_/Q vssd1 vssd1 vccd1 vccd1 _3430_/A sky130_fd_sc_hd__xnor2_2
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4965_ _4955_/X _4968_/C _4968_/B vssd1 vssd1 vccd1 vccd1 _4966_/C sky130_fd_sc_hd__a21oi_1
XFILLER_51_234 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3916_ _3872_/X _3874_/X _3917_/A vssd1 vssd1 vccd1 vccd1 _3916_/X sky130_fd_sc_hd__a21o_1
XFILLER_51_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4343__A _4397_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4896_ _5983_/Q _4854_/X _4855_/X vssd1 vssd1 vccd1 vccd1 _4896_/X sky130_fd_sc_hd__o21a_1
XFILLER_32_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3847_ _4556_/B _4474_/C vssd1 vssd1 vccd1 vccd1 _5261_/A sky130_fd_sc_hd__nand2_1
XFILLER_22_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3778_ _3784_/A _3778_/B vssd1 vssd1 vccd1 vccd1 _3779_/A sky130_fd_sc_hd__and2_1
X_5517_ _6073_/Q _5526_/B vssd1 vssd1 vccd1 vccd1 _5517_/X sky130_fd_sc_hd__or2_1
XANTENNA__5174__A _5174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5448_ _5579_/A _5469_/B vssd1 vssd1 vccd1 vccd1 _5449_/A sky130_fd_sc_hd__or2_1
X_5379_ _5579_/A _5379_/B vssd1 vssd1 vccd1 vccd1 _5399_/B sky130_fd_sc_hd__nor2_1
XFILLER_59_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4456__C1 _3269_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4223__A2 _3938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5349__A _5405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4399__S _4399_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4750_ _6103_/Q _4749_/X _4771_/S vssd1 vssd1 vccd1 vccd1 _4750_/X sky130_fd_sc_hd__mux2_1
X_3701_ _3701_/A _3701_/B vssd1 vssd1 vccd1 vccd1 _3702_/A sky130_fd_sc_hd__and2_1
X_4681_ _4781_/A vssd1 vssd1 vccd1 vccd1 _4720_/S sky130_fd_sc_hd__clkbuf_2
X_3632_ _3632_/A _3632_/B vssd1 vssd1 vccd1 vccd1 _3633_/A sky130_fd_sc_hd__and2_1
X_5302_ _2931_/B _3486_/A _5301_/X _5299_/Y vssd1 vssd1 vccd1 vccd1 _5302_/X sky130_fd_sc_hd__o211a_1
XANTENNA__4102__S _4116_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3563_ _3563_/A vssd1 vssd1 vccd1 vccd1 _3563_/X sky130_fd_sc_hd__buf_2
X_3494_ _3494_/A _3494_/B vssd1 vssd1 vccd1 vccd1 _3494_/Y sky130_fd_sc_hd__nor2_1
XFILLER_5_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5233_ _5233_/A _5233_/B _5233_/C _3861_/A vssd1 vssd1 vccd1 vccd1 _5236_/C sky130_fd_sc_hd__or4b_1
XFILLER_68_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5164_ _5984_/Q _5168_/B vssd1 vssd1 vccd1 vccd1 _5164_/X sky130_fd_sc_hd__or2_1
XFILLER_68_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4115_ _6114_/Q _5776_/Q _4128_/S vssd1 vssd1 vccd1 vccd1 _4115_/X sky130_fd_sc_hd__mux2_1
X_5095_ _5960_/Q _5100_/B vssd1 vssd1 vccd1 vccd1 _5095_/X sky130_fd_sc_hd__or2_1
XFILLER_83_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4046_ _5757_/Q _4045_/X _4046_/S vssd1 vssd1 vccd1 vccd1 _4047_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5997_ _6002_/CLK _5997_/D vssd1 vssd1 vccd1 vccd1 _5997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5402__A1 _3582_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5169__A _5391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4948_ _4948_/A vssd1 vssd1 vccd1 vccd1 _4948_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_12_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4879_ _5903_/Q _4858_/X _4877_/X _4878_/X vssd1 vssd1 vccd1 vccd1 _5903_/D sky130_fd_sc_hd__a22o_1
XFILLER_58_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2975__B _4218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_10 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5079__A _5601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_proj_example_201 vssd1 vssd1 vccd1 vccd1 user_proj_example_201/HI la_data_out[108]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_212 vssd1 vssd1 vccd1 vccd1 user_proj_example_212/HI la_data_out[119]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_245 vssd1 vssd1 vccd1 vccd1 user_proj_example_245/HI wbs_dat_o[24]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_234 vssd1 vssd1 vccd1 vccd1 user_proj_example_234/HI wbs_dat_o[13]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_223 vssd1 vssd1 vccd1 vccd1 user_proj_example_223/HI wbs_dat_o[2]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_278 vssd1 vssd1 vccd1 vccd1 io_out[26] user_proj_example_278/LO
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_267 vssd1 vssd1 vccd1 vccd1 io_out[15] user_proj_example_267/LO
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_256 vssd1 vssd1 vccd1 vccd1 io_out[4] user_proj_example_256/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA__4904__B1 _4607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5920_ _5920_/CLK _5920_/D vssd1 vssd1 vccd1 vccd1 _5920_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5632__A1 _5357_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5851_ _6005_/CLK _5851_/D vssd1 vssd1 vccd1 vccd1 _5851_/Q sky130_fd_sc_hd__dfxtp_1
X_2994_ _3049_/A _2994_/B vssd1 vssd1 vccd1 vccd1 _3845_/C sky130_fd_sc_hd__nand2_1
X_5782_ _6005_/CLK _5782_/D vssd1 vssd1 vccd1 vccd1 _5782_/Q sky130_fd_sc_hd__dfxtp_1
X_4802_ _6060_/Q _4757_/X _4767_/X _4801_/X vssd1 vssd1 vccd1 vccd1 _4802_/X sky130_fd_sc_hd__a211o_1
XFILLER_21_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4733_ _4717_/X _4731_/X _4732_/X _4722_/X vssd1 vssd1 vccd1 vccd1 _4733_/X sky130_fd_sc_hd__o211a_1
X_4664_ _4716_/A vssd1 vssd1 vccd1 vccd1 _4664_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4595_ _4842_/A vssd1 vssd1 vccd1 vccd1 _4917_/B sky130_fd_sc_hd__clkbuf_2
X_3615_ _5664_/Q _3618_/B vssd1 vssd1 vccd1 vccd1 _3615_/X sky130_fd_sc_hd__or2_1
X_3546_ _3546_/A vssd1 vssd1 vccd1 vccd1 _3546_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3477_ _3820_/B _2969_/B _3476_/X _4229_/A vssd1 vssd1 vccd1 vccd1 _3477_/X sky130_fd_sc_hd__a31o_1
X_5216_ _5065_/A _6001_/Q _5216_/S vssd1 vssd1 vccd1 vccd1 _5217_/B sky130_fd_sc_hd__mux2_1
XFILLER_69_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5147_ _5345_/A vssd1 vssd1 vccd1 vccd1 _5405_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_28_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5078_ _5603_/B vssd1 vssd1 vccd1 vccd1 _5601_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_71_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4029_ _4029_/A vssd1 vssd1 vccd1 vccd1 _5752_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5627__A _5638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2986__A _3049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input34_A la_data_in[59] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4706__A _4706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3400_ _5277_/A _3400_/B _2846_/C vssd1 vssd1 vccd1 vccd1 _3502_/A sky130_fd_sc_hd__or3b_2
X_4380_ _6052_/Q _5829_/Q _4380_/S vssd1 vssd1 vccd1 vccd1 _4380_/X sky130_fd_sc_hd__mux2_1
X_3331_ _4113_/A vssd1 vssd1 vccd1 vccd1 _3331_/X sky130_fd_sc_hd__clkbuf_2
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ _3374_/A vssd1 vssd1 vccd1 vccd1 _3509_/A sky130_fd_sc_hd__clkbuf_2
X_6050_ _6050_/CLK _6050_/D vssd1 vssd1 vccd1 vccd1 _6050_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3193_ _5921_/Q _5912_/Q vssd1 vssd1 vccd1 vccd1 _3193_/X sky130_fd_sc_hd__xor2_1
X_5001_ _5932_/Q _4999_/A _4990_/X vssd1 vssd1 vccd1 vccd1 _5002_/B sky130_fd_sc_hd__o21ai_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4616__A _4842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5903_ _5983_/CLK _5903_/D vssd1 vssd1 vccd1 vccd1 _5903_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5834_ _6050_/CLK _5834_/D vssd1 vssd1 vccd1 vccd1 _5834_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4041__A0 _6098_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2977_ _5848_/Q vssd1 vssd1 vccd1 vccd1 _3873_/A sky130_fd_sc_hd__clkinv_2
X_5765_ _6109_/CLK _5765_/D vssd1 vssd1 vccd1 vccd1 _5765_/Q sky130_fd_sc_hd__dfxtp_1
X_4716_ _4716_/A vssd1 vssd1 vccd1 vccd1 _4716_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5696_ _6031_/CLK _5696_/D vssd1 vssd1 vccd1 vccd1 _5696_/Q sky130_fd_sc_hd__dfxtp_1
X_4647_ _6093_/Q _4646_/X _4668_/S vssd1 vssd1 vccd1 vccd1 _4647_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4578_ _4858_/A vssd1 vssd1 vccd1 vccd1 _4756_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3529_ _3529_/A _3529_/B vssd1 vssd1 vccd1 vccd1 _3529_/Y sky130_fd_sc_hd__nor2_1
XFILLER_1_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_27_wb_clk_i clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5920_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_40_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5357__A input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4335__B2 _6066_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3543__C1 _3408_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4099__A0 _5959_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4200__S _4200_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4436__A _4436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2882__C _3256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_340 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2900_ _2885_/Y _2892_/X _3158_/A vssd1 vssd1 vccd1 vccd1 _2900_/Y sky130_fd_sc_hd__o21ai_1
X_3880_ _3878_/X _3879_/Y _3880_/S vssd1 vssd1 vccd1 vccd1 _3880_/X sky130_fd_sc_hd__mux2_1
X_2831_ _3117_/A vssd1 vssd1 vccd1 vccd1 _3272_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5550_ _3607_/X _5536_/X _5549_/X _5545_/X vssd1 vssd1 vccd1 vccd1 _6085_/D sky130_fd_sc_hd__o211a_1
X_4501_ _5744_/Q _4501_/B _5737_/Q _4500_/Y vssd1 vssd1 vccd1 vccd1 _4502_/C sky130_fd_sc_hd__or4b_1
X_5481_ _6060_/Q _5483_/B vssd1 vssd1 vccd1 vccd1 _5481_/X sky130_fd_sc_hd__or2_1
X_4432_ _5975_/Q _5845_/Q _4432_/S vssd1 vssd1 vccd1 vccd1 _4432_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4363_ _6047_/Q _5824_/Q _4363_/S vssd1 vssd1 vccd1 vccd1 _4363_/X sky130_fd_sc_hd__mux2_1
X_3314_ _3427_/C _3483_/B _3843_/B vssd1 vssd1 vccd1 vccd1 _3314_/X sky130_fd_sc_hd__a21o_1
X_4294_ _4294_/A _4294_/B _4294_/C _4294_/D vssd1 vssd1 vccd1 vccd1 _4294_/X sky130_fd_sc_hd__and4_1
XANTENNA__4110__S _4110_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6102_ _6135_/CLK _6102_/D vssd1 vssd1 vccd1 vccd1 _6102_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3245_ _3632_/A vssd1 vssd1 vccd1 vccd1 _3245_/X sky130_fd_sc_hd__clkbuf_2
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6033_ _6108_/CLK _6033_/D vssd1 vssd1 vccd1 vccd1 _6033_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3176_ _5913_/Q vssd1 vssd1 vccd1 vccd1 _4935_/A sky130_fd_sc_hd__inv_2
XFILLER_54_424 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5817_ _6005_/CLK _5817_/D vssd1 vssd1 vccd1 vccd1 _5817_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5177__A _5186_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4565__A1 _3135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5748_ _5796_/CLK _5748_/D vssd1 vssd1 vccd1 vccd1 _5748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4317__A1 _3494_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5679_ _5703_/CLK _5679_/D vssd1 vssd1 vccd1 vccd1 _5679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5640__A _6119_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4005__B1 _4452_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput70 _5897_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[84] sky130_fd_sc_hd__buf_2
Xoutput81 _5908_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[95] sky130_fd_sc_hd__buf_2
XFILLER_68_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4492__B1 _5171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3030_ _3264_/A _3035_/C vssd1 vssd1 vccd1 vccd1 _3037_/B sky130_fd_sc_hd__nand2_1
XFILLER_48_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_3_0__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4981_ _5011_/A _4981_/B vssd1 vssd1 vccd1 vccd1 _4995_/B sky130_fd_sc_hd__nor2_2
XFILLER_23_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3932_ _3932_/A vssd1 vssd1 vccd1 vccd1 _3932_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4795__A1 _6035_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3863_ _5233_/A _4010_/A _3902_/B vssd1 vssd1 vccd1 vccd1 _3888_/A sky130_fd_sc_hd__or3_1
XANTENNA__4105__S _4116_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5602_ _5602_/A vssd1 vssd1 vccd1 vccd1 _5602_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3794_ _3794_/A vssd1 vssd1 vccd1 vccd1 _5171_/B sky130_fd_sc_hd__inv_2
X_5533_ _6080_/Q _5533_/B vssd1 vssd1 vccd1 vccd1 _5533_/X sky130_fd_sc_hd__or2_1
X_5464_ _5396_/X _5449_/A _5463_/X _5461_/X vssd1 vssd1 vccd1 vccd1 _6054_/D sky130_fd_sc_hd__o211a_1
X_5395_ _5393_/X _5378_/X _5394_/X _5391_/X vssd1 vssd1 vccd1 vccd1 _6029_/D sky130_fd_sc_hd__o211a_1
X_4415_ _4415_/A vssd1 vssd1 vccd1 vccd1 _5840_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3245__A _3632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4346_ _6042_/Q _5819_/Q _5278_/A vssd1 vssd1 vccd1 vccd1 _4346_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4277_ _5736_/Q vssd1 vssd1 vccd1 vccd1 _4277_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4483__B1 _3245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6016_ _6018_/CLK _6016_/D vssd1 vssd1 vccd1 vccd1 _6016_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3228_ _6034_/Q _5935_/Q vssd1 vssd1 vccd1 vccd1 _3228_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_82_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3159_ _3873_/A _3159_/B vssd1 vssd1 vccd1 vccd1 _3257_/A sky130_fd_sc_hd__nor2_1
XFILLER_27_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4786__A1 _6034_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4804__A _4855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5499__C1 _5488_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3155__A _4251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_59_wb_clk_i_A clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2994__A _3049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5370__A _6023_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3277__A1 _4220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_42_wb_clk_i clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5999_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4226__B1 _4452_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5423__C1 _5420_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3201__B2 _5354_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3201__A1 _6023_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5545__A _5597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4200_ _5802_/Q _4199_/X _4200_/S vssd1 vssd1 vccd1 vccd1 _4201_/A sky130_fd_sc_hd__mux2_1
X_5180_ _5186_/A _5180_/B vssd1 vssd1 vccd1 vccd1 _5181_/A sky130_fd_sc_hd__and2_1
XFILLER_3_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4131_ _4182_/A vssd1 vssd1 vccd1 vccd1 _4145_/S sky130_fd_sc_hd__clkbuf_2
X_4062_ _6105_/Q _3869_/A _4075_/S vssd1 vssd1 vccd1 vccd1 _4062_/X sky130_fd_sc_hd__mux2_1
X_3013_ _3841_/A _3839_/B vssd1 vssd1 vccd1 vccd1 _3428_/B sky130_fd_sc_hd__xnor2_2
XFILLER_64_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4964_ _4968_/B _4964_/B _4968_/C vssd1 vssd1 vccd1 vccd1 _4966_/B sky130_fd_sc_hd__and3_1
XFILLER_51_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3915_ _3915_/A vssd1 vssd1 vccd1 vccd1 _5720_/D sky130_fd_sc_hd__clkbuf_1
X_4895_ _5975_/Q _4859_/X _4869_/X _4894_/X vssd1 vssd1 vccd1 vccd1 _4895_/X sky130_fd_sc_hd__a211o_1
X_3846_ _4283_/A _4471_/A _4283_/B _4283_/C _3845_/X vssd1 vssd1 vccd1 vccd1 _4474_/C
+ sky130_fd_sc_hd__o41a_1
X_3777_ _3604_/A _5708_/Q _3780_/S vssd1 vssd1 vccd1 vccd1 _3778_/B sky130_fd_sc_hd__mux2_1
X_5516_ _5533_/B vssd1 vssd1 vccd1 vccd1 _5526_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__5174__B _5201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5447_ _5373_/X _5427_/A _5445_/X _5446_/X vssd1 vssd1 vccd1 vccd1 _6048_/D sky130_fd_sc_hd__o211a_1
XFILLER_59_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5378_ _5401_/B vssd1 vssd1 vccd1 vccd1 _5378_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4329_ _4555_/B _4329_/B vssd1 vssd1 vccd1 vccd1 _4329_/Y sky130_fd_sc_hd__nor2_1
XFILLER_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5653__C1 _5172_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3700_ _3611_/A _5687_/Q _3707_/S vssd1 vssd1 vccd1 vccd1 _3701_/B sky130_fd_sc_hd__mux2_1
X_4680_ _6120_/Q _4678_/X _4719_/S vssd1 vssd1 vccd1 vccd1 _4680_/X sky130_fd_sc_hd__mux2_1
X_3631_ input6/X _5667_/Q _3641_/S vssd1 vssd1 vccd1 vccd1 _3632_/B sky130_fd_sc_hd__mux2_1
X_3562_ _5744_/Q _3412_/X _3561_/Y _3255_/X vssd1 vssd1 vccd1 vccd1 _5744_/D sky130_fd_sc_hd__a22o_1
X_5301_ _5301_/A _5301_/B _5301_/C vssd1 vssd1 vccd1 vccd1 _5301_/X sky130_fd_sc_hd__and3_1
X_3493_ _3493_/A vssd1 vssd1 vccd1 vccd1 _3493_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5232_ _5657_/Q _3061_/A _5231_/X vssd1 vssd1 vccd1 vccd1 _5232_/X sky130_fd_sc_hd__a21o_1
XFILLER_68_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5163_ _5065_/X _5149_/X _5162_/X _5158_/X vssd1 vssd1 vccd1 vccd1 _5983_/D sky130_fd_sc_hd__o211a_1
XFILLER_68_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4114_ _4182_/A vssd1 vssd1 vccd1 vccd1 _4128_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_56_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5094_ _5065_/X _5080_/X _5093_/X _5087_/X vssd1 vssd1 vccd1 vccd1 _5959_/D sky130_fd_sc_hd__o211a_1
X_4045_ _6099_/Q _5756_/Q _4058_/S vssd1 vssd1 vccd1 vccd1 _4045_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5996_ _5996_/CLK _5996_/D vssd1 vssd1 vccd1 vccd1 _5996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3413__A1 _3391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4947_ _4954_/A _4972_/B vssd1 vssd1 vccd1 vccd1 _4948_/A sky130_fd_sc_hd__nor2_1
X_4878_ _5981_/Q _4854_/X _4855_/X vssd1 vssd1 vccd1 vccd1 _4878_/X sky130_fd_sc_hd__o21a_1
X_3829_ _4281_/A _5719_/Q _4283_/B _3829_/D vssd1 vssd1 vccd1 vccd1 _3830_/B sky130_fd_sc_hd__or4_1
XFILLER_20_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_proj_example_202 vssd1 vssd1 vccd1 vccd1 user_proj_example_202/HI la_data_out[109]
+ sky130_fd_sc_hd__conb_1
XANTENNA__4203__S _4203_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xuser_proj_example_213 vssd1 vssd1 vccd1 vccd1 user_proj_example_213/HI la_data_out[120]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_224 vssd1 vssd1 vccd1 vccd1 user_proj_example_224/HI wbs_dat_o[3]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_246 vssd1 vssd1 vccd1 vccd1 user_proj_example_246/HI wbs_dat_o[25]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_235 vssd1 vssd1 vccd1 vccd1 user_proj_example_235/HI wbs_dat_o[14]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_279 vssd1 vssd1 vccd1 vccd1 io_out[27] user_proj_example_279/LO
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_268 vssd1 vssd1 vccd1 vccd1 io_out[16] user_proj_example_268/LO
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_257 vssd1 vssd1 vccd1 vccd1 io_out[5] user_proj_example_257/LO
+ sky130_fd_sc_hd__conb_1
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3340__B1 _5258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4840__A0 _5665_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5850_ _6131_/CLK _5850_/D vssd1 vssd1 vccd1 vccd1 _5850_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2993_ _3005_/C vssd1 vssd1 vccd1 vccd1 _3484_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_396 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4801_ _4768_/X _4799_/X _4800_/X _4773_/X vssd1 vssd1 vccd1 vccd1 _4801_/X sky130_fd_sc_hd__o211a_1
X_5781_ _6117_/CLK _5781_/D vssd1 vssd1 vccd1 vccd1 _5781_/Q sky130_fd_sc_hd__dfxtp_1
X_4732_ _6077_/Q _4732_/B vssd1 vssd1 vccd1 vccd1 _4732_/X sky130_fd_sc_hd__or2_1
X_4663_ _5882_/Q _4653_/X _4661_/X _4662_/X vssd1 vssd1 vccd1 vccd1 _5882_/D sky130_fd_sc_hd__a22o_1
XANTENNA__3518__A _3518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3614_ _3614_/A vssd1 vssd1 vccd1 vccd1 _3614_/X sky130_fd_sc_hd__clkbuf_2
X_4594_ _4594_/A _4594_/B _4594_/C vssd1 vssd1 vccd1 vccd1 _4842_/A sky130_fd_sc_hd__or3_2
X_3545_ _3221_/X _3532_/X _3544_/X vssd1 vssd1 vccd1 vccd1 _5739_/D sky130_fd_sc_hd__a21bo_1
X_3476_ _5279_/A _3824_/D _3476_/C _3282_/A vssd1 vssd1 vccd1 vccd1 _3476_/X sky130_fd_sc_hd__or4b_1
X_5215_ _5215_/A vssd1 vssd1 vccd1 vccd1 _6000_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4349__A _4366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3882__A1 _3867_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5146_ _5075_/X _5125_/A _5145_/X _5141_/X vssd1 vssd1 vccd1 vccd1 _5978_/D sky130_fd_sc_hd__o211a_1
XFILLER_28_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5608__C1 _5597_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3882__B2 _5761_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5077_ _5075_/X _5050_/A _5076_/X _5067_/X vssd1 vssd1 vccd1 vccd1 _5954_/D sky130_fd_sc_hd__o211a_1
XFILLER_84_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4028_ _5752_/Q _4027_/X _4028_/S vssd1 vssd1 vccd1 vccd1 _4029_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5979_ _5983_/CLK _5979_/D vssd1 vssd1 vccd1 vccd1 _5979_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_536 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4259__A _4259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input27_A la_data_in[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4722__A _4824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5537__B _5537_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3330_ _4287_/A vssd1 vssd1 vccd1 vccd1 _4113_/A sky130_fd_sc_hd__clkbuf_2
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3261_ _3522_/B _3260_/X _3117_/Y _3423_/C vssd1 vssd1 vccd1 vccd1 _3261_/X sky130_fd_sc_hd__a22o_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _5932_/Q _5931_/Q _5000_/C vssd1 vssd1 vccd1 vccd1 _5006_/C sky130_fd_sc_hd__and3_1
XFILLER_85_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3192_ _5918_/Q _5909_/Q vssd1 vssd1 vccd1 vccd1 _3192_/X sky130_fd_sc_hd__or2_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3616__A1 _3614_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4108__S _4116_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5902_ _5983_/CLK _5902_/D vssd1 vssd1 vccd1 vccd1 _5902_/Q sky130_fd_sc_hd__dfxtp_1
X_5833_ _6050_/CLK _5833_/D vssd1 vssd1 vccd1 vccd1 _5833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2976_ _5718_/Q vssd1 vssd1 vccd1 vccd1 _4217_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5764_ _6109_/CLK _5764_/D vssd1 vssd1 vccd1 vccd1 _5764_/Q sky130_fd_sc_hd__dfxtp_1
X_4715_ _5887_/Q _4705_/X _4713_/X _4714_/Y vssd1 vssd1 vccd1 vccd1 _5887_/D sky130_fd_sc_hd__a22o_1
X_5695_ _6027_/CLK _5695_/D vssd1 vssd1 vccd1 vccd1 _5695_/Q sky130_fd_sc_hd__dfxtp_1
X_4646_ _6117_/Q _4645_/X _4667_/S vssd1 vssd1 vccd1 vccd1 _4646_/X sky130_fd_sc_hd__mux2_1
X_4577_ input3/X _4577_/B input2/X _3564_/B vssd1 vssd1 vccd1 vccd1 _4858_/A sky130_fd_sc_hd__or4b_4
XANTENNA__3552__B1 _3245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5463__A _6054_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3528_ _5862_/Q _5861_/Q _5860_/Q _5863_/Q vssd1 vssd1 vccd1 vccd1 _3529_/B sky130_fd_sc_hd__or4bb_1
X_3459_ _5279_/A _3482_/A _3841_/B _3459_/D vssd1 vssd1 vccd1 vccd1 _3460_/D sky130_fd_sc_hd__or4_1
XFILLER_69_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5129_ _5971_/Q _5138_/B vssd1 vssd1 vccd1 vccd1 _5129_/X sky130_fd_sc_hd__or2_1
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4807__A _4858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5638__A _5638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5532__A1 _3563_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5373__A _5373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4717__A _4717_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2830_ _3929_/B _5245_/A vssd1 vssd1 vccd1 vccd1 _3117_/A sky130_fd_sc_hd__nand2_1
XFILLER_16_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4500_ _4496_/Y _5738_/Q _3553_/X vssd1 vssd1 vccd1 vccd1 _4500_/Y sky130_fd_sc_hd__a21oi_1
X_5480_ _3601_/X _5470_/X _5479_/X _5477_/X vssd1 vssd1 vccd1 vccd1 _6059_/D sky130_fd_sc_hd__o211a_1
XANTENNA__4326__A2 _3484_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4431_ _4431_/A vssd1 vssd1 vccd1 vccd1 _5845_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5523__A1 _5386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4362_ _4362_/A vssd1 vssd1 vccd1 vccd1 _5824_/D sky130_fd_sc_hd__clkbuf_1
X_3313_ _3326_/A _3430_/A vssd1 vssd1 vccd1 vccd1 _3843_/B sky130_fd_sc_hd__and2_1
X_4293_ _4293_/A _4327_/A vssd1 vssd1 vccd1 vccd1 _4294_/D sky130_fd_sc_hd__or2_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6101_ _6101_/CLK _6101_/D vssd1 vssd1 vccd1 vccd1 _6101_/Q sky130_fd_sc_hd__dfxtp_1
X_3244_ _4982_/B _4954_/A _3244_/C vssd1 vssd1 vccd1 vccd1 _4981_/B sky130_fd_sc_hd__and3_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6032_ _6040_/CLK _6032_/D vssd1 vssd1 vccd1 vccd1 _6032_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3175_ _5922_/Q vssd1 vssd1 vccd1 vccd1 _4968_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5816_ _6005_/CLK _5816_/D vssd1 vssd1 vccd1 vccd1 _5816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5747_ _6121_/CLK _5747_/D vssd1 vssd1 vccd1 vccd1 _5747_/Q sky130_fd_sc_hd__dfxtp_1
X_2959_ _3044_/D _3322_/A _2959_/C _4464_/B vssd1 vssd1 vccd1 vccd1 _3283_/B sky130_fd_sc_hd__nor4_4
XFILLER_22_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5678_ _5703_/CLK _5678_/D vssd1 vssd1 vccd1 vccd1 _5678_/Q sky130_fd_sc_hd__dfxtp_1
X_4629_ _4781_/A vssd1 vssd1 vccd1 vccd1 _4668_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_89_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_49_wb_clk_i_A clkbuf_3_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_49_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3798__D _4607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4272__A _4970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3335__B _5258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput60 _5887_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[74] sky130_fd_sc_hd__buf_2
XFILLER_68_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput71 _5898_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[85] sky130_fd_sc_hd__buf_2
Xoutput82 _5987_/Q vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__buf_2
XANTENNA__3819__A1 _5336_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output58_A _5885_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4980_ _3180_/Y _4972_/B _4976_/Y _4979_/X _3255_/X vssd1 vssd1 vccd1 vccd1 _5926_/D
+ sky130_fd_sc_hd__o311a_1
X_3931_ _3964_/A vssd1 vssd1 vccd1 vccd1 _3932_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__5278__A _5278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3862_ _3484_/B _4220_/B _5234_/B _3861_/X vssd1 vssd1 vccd1 vccd1 _3902_/B sky130_fd_sc_hd__o31ai_1
XANTENNA__4182__A _4182_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5601_ _5601_/A _5601_/B vssd1 vssd1 vccd1 vccd1 _5602_/A sky130_fd_sc_hd__or2_1
XFILLER_31_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3793_ _3793_/A vssd1 vssd1 vccd1 vccd1 _5712_/D sky130_fd_sc_hd__clkbuf_1
X_5532_ _3563_/X _5514_/A _5531_/X _5529_/X vssd1 vssd1 vccd1 vccd1 _6079_/D sky130_fd_sc_hd__o211a_1
X_5463_ _6054_/Q _5467_/B vssd1 vssd1 vccd1 vccd1 _5463_/X sky130_fd_sc_hd__or2_1
X_5394_ _6029_/Q _5399_/B vssd1 vssd1 vccd1 vccd1 _5394_/X sky130_fd_sc_hd__or2_1
X_4414_ _5840_/Q _4413_/X _4417_/S vssd1 vssd1 vccd1 vccd1 _4415_/A sky130_fd_sc_hd__mux2_1
X_4345_ _4345_/A vssd1 vssd1 vccd1 vccd1 _5819_/D sky130_fd_sc_hd__clkbuf_1
X_4276_ _4276_/A _4276_/B _4276_/C vssd1 vssd1 vccd1 vccd1 _5808_/D sky130_fd_sc_hd__nor3_1
X_6015_ _6018_/CLK _6015_/D vssd1 vssd1 vccd1 vccd1 _6015_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3227_ _6027_/Q vssd1 vssd1 vccd1 vccd1 _5387_/A sky130_fd_sc_hd__clkinv_2
XFILLER_39_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3158_ _3158_/A vssd1 vssd1 vccd1 vccd1 _3522_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_54_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3089_ _4237_/C vssd1 vssd1 vccd1 vccd1 _3423_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5188__A _5188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_5_wb_clk_i_A clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_2_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2994__B _2994_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3277__A2 _3275_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_11_wb_clk_i _5813_/CLK vssd1 vssd1 vccd1 vccd1 _5736_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4130_ _4130_/A vssd1 vssd1 vccd1 vccd1 _5781_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3081__A _3480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4061_ _4095_/A vssd1 vssd1 vccd1 vccd1 _4075_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_3_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3012_ _3838_/A _5228_/B _3288_/C vssd1 vssd1 vccd1 vccd1 _3841_/C sky130_fd_sc_hd__or3_2
XFILLER_76_391 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4963_ _4966_/A _4963_/B vssd1 vssd1 vccd1 vccd1 _5921_/D sky130_fd_sc_hd__nor2_1
XFILLER_36_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3914_ _3910_/X _3897_/B _3914_/S vssd1 vssd1 vccd1 vccd1 _3915_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4116__S _4116_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4894_ _4870_/X _4892_/X _4893_/X _4875_/X vssd1 vssd1 vccd1 vccd1 _4894_/X sky130_fd_sc_hd__o211a_1
X_3845_ _3845_/A _4438_/B _3845_/C _3845_/D vssd1 vssd1 vccd1 vccd1 _3845_/X sky130_fd_sc_hd__or4_1
XANTENNA__3728__A0 _5366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3776_ _3776_/A vssd1 vssd1 vccd1 vccd1 _5707_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4640__A _6068_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5515_ _5581_/A _5535_/B vssd1 vssd1 vccd1 vccd1 _5533_/B sky130_fd_sc_hd__nor2_1
XANTENNA__3256__A _3256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5446_ _5461_/A vssd1 vssd1 vccd1 vccd1 _5446_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5377_ _5581_/A _5405_/B vssd1 vssd1 vccd1 vccd1 _5401_/B sky130_fd_sc_hd__or2_1
XFILLER_86_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4328_ _3929_/C _4327_/A _4319_/X _4325_/X _4327_/Y vssd1 vssd1 vccd1 vccd1 _4328_/X
+ sky130_fd_sc_hd__a41o_1
XANTENNA_input1_A io_in[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4259_ _4259_/A _4259_/B vssd1 vssd1 vccd1 vccd1 _4259_/Y sky130_fd_sc_hd__nor2_1
XFILLER_74_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4456__A1 _3469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3719__A0 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3166__A _3553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4695__A1 _6025_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5556__A _5597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3630_ _3630_/A vssd1 vssd1 vccd1 vccd1 _5666_/D sky130_fd_sc_hd__clkbuf_1
X_3561_ _3561_/A _3561_/B vssd1 vssd1 vccd1 vccd1 _3561_/Y sky130_fd_sc_hd__nor2_1
X_5300_ _5269_/B _5278_/B _5257_/B _5299_/Y vssd1 vssd1 vccd1 vccd1 _5307_/A sky130_fd_sc_hd__o31a_1
XFILLER_52_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3492_ _3505_/C _3425_/X _3489_/X _3491_/X vssd1 vssd1 vccd1 vccd1 _6122_/D sky130_fd_sc_hd__a22o_1
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5231_ _5789_/Q _5229_/Y _5230_/X _3331_/X vssd1 vssd1 vccd1 vccd1 _5231_/X sky130_fd_sc_hd__o211a_1
XANTENNA__4686__A1 _6024_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5162_ _5983_/Q _5162_/B vssd1 vssd1 vccd1 vccd1 _5162_/X sky130_fd_sc_hd__or2_1
X_4113_ _4113_/A vssd1 vssd1 vccd1 vccd1 _4182_/A sky130_fd_sc_hd__buf_2
X_5093_ _5959_/Q _5093_/B vssd1 vssd1 vccd1 vccd1 _5093_/X sky130_fd_sc_hd__or2_1
XFILLER_83_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4044_ _4095_/A vssd1 vssd1 vccd1 vccd1 _4058_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_49_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5995_ _6003_/CLK _5995_/D vssd1 vssd1 vccd1 vccd1 _5995_/Q sky130_fd_sc_hd__dfxtp_1
X_4946_ _5855_/Q _5854_/Q _4946_/C vssd1 vssd1 vccd1 vccd1 _4972_/B sky130_fd_sc_hd__nor3_2
XFILLER_33_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4877_ _5973_/Q _4859_/X _4869_/X _4876_/X vssd1 vssd1 vccd1 vccd1 _4877_/X sky130_fd_sc_hd__a211o_1
X_3828_ _2982_/B _3828_/B _4470_/B _5247_/B vssd1 vssd1 vccd1 vccd1 _5233_/B sky130_fd_sc_hd__and4b_1
XFILLER_20_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3759_ _3563_/A _5703_/Q _3762_/S vssd1 vssd1 vccd1 vccd1 _3760_/B sky130_fd_sc_hd__mux2_1
XANTENNA__4913__A2 _4623_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4677__A1 _5883_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5429_ _5445_/B vssd1 vssd1 vccd1 vccd1 _5439_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__3714__A _5343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_180 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_proj_example_203 vssd1 vssd1 vccd1 vccd1 user_proj_example_203/HI la_data_out[110]
+ sky130_fd_sc_hd__conb_1
XFILLER_23_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_proj_example_236 vssd1 vssd1 vccd1 vccd1 user_proj_example_236/HI wbs_dat_o[15]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_225 vssd1 vssd1 vccd1 vccd1 user_proj_example_225/HI wbs_dat_o[4]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_214 vssd1 vssd1 vccd1 vccd1 user_proj_example_214/HI la_data_out[121]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_269 vssd1 vssd1 vccd1 vccd1 io_out[17] user_proj_example_269/LO
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_258 vssd1 vssd1 vccd1 vccd1 io_out[6] user_proj_example_258/LO
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_247 vssd1 vssd1 vccd1 vccd1 user_proj_example_247/HI wbs_dat_o[26]
+ sky130_fd_sc_hd__conb_1
XANTENNA__4904__A2 _5379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3340__A1 _4220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4800_ _6084_/Q _4834_/B vssd1 vssd1 vccd1 vccd1 _4800_/X sky130_fd_sc_hd__or2_1
X_2992_ _3256_/A _3296_/B vssd1 vssd1 vccd1 vccd1 _3005_/C sky130_fd_sc_hd__nand2_1
XFILLER_61_364 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5780_ _6117_/CLK _5780_/D vssd1 vssd1 vccd1 vccd1 _5780_/Q sky130_fd_sc_hd__dfxtp_1
X_4731_ _6101_/Q _4729_/X _4771_/S vssd1 vssd1 vccd1 vccd1 _4731_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4662_ _6022_/Q _4606_/X _4607_/X vssd1 vssd1 vccd1 vccd1 _4662_/X sky130_fd_sc_hd__o21a_1
X_3613_ _3611_/X _3592_/A _3612_/X _3609_/X vssd1 vssd1 vccd1 vccd1 _5663_/D sky130_fd_sc_hd__o211a_1
X_4593_ _6089_/Q _4590_/X _4781_/A vssd1 vssd1 vccd1 vccd1 _4593_/X sky130_fd_sc_hd__mux2_1
X_3544_ _4567_/A _3544_/B _3544_/C _3544_/D vssd1 vssd1 vccd1 vccd1 _3544_/X sky130_fd_sc_hd__or4_1
XANTENNA__4108__A0 _5775_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5305__C1 _3867_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3475_ _3435_/A _3440_/B _3474_/X _3480_/C vssd1 vssd1 vccd1 vccd1 _3475_/X sky130_fd_sc_hd__o22a_1
X_5214_ _5220_/A _5214_/B vssd1 vssd1 vccd1 vccd1 _5215_/A sky130_fd_sc_hd__and2_1
XFILLER_69_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5145_ _5978_/Q _5145_/B vssd1 vssd1 vccd1 vccd1 _5145_/X sky130_fd_sc_hd__or2_1
XFILLER_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5076_ _5954_/Q _5076_/B vssd1 vssd1 vccd1 vccd1 _5076_/X sky130_fd_sc_hd__or2_1
XANTENNA__5084__A1 _5045_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4027_ _6093_/Q _4014_/X _5751_/Q _4017_/X vssd1 vssd1 vccd1 vccd1 _4027_/X sky130_fd_sc_hd__a22o_1
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5978_ _5986_/CLK _5978_/D vssd1 vssd1 vccd1 vccd1 _5978_/Q sky130_fd_sc_hd__dfxtp_1
X_4929_ _5067_/A vssd1 vssd1 vccd1 vccd1 _4929_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_12_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3354__A _3897_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ _4322_/B vssd1 vssd1 vccd1 vccd1 _3260_/X sky130_fd_sc_hd__clkbuf_2
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3191_ _5918_/Q _5909_/Q vssd1 vssd1 vccd1 vccd1 _3191_/Y sky130_fd_sc_hd__nand2_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5901_ _5966_/CLK _5901_/D vssd1 vssd1 vccd1 vccd1 _5901_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_331 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5832_ _6050_/CLK _5832_/D vssd1 vssd1 vccd1 vccd1 _5832_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5763_ _6109_/CLK _5763_/D vssd1 vssd1 vccd1 vccd1 _5763_/Q sky130_fd_sc_hd__dfxtp_1
X_2975_ _3826_/C _4218_/B vssd1 vssd1 vccd1 vccd1 _2975_/Y sky130_fd_sc_hd__nand2_1
X_4714_ _5387_/A _4602_/X _4623_/X vssd1 vssd1 vccd1 vccd1 _4714_/Y sky130_fd_sc_hd__a21oi_1
X_5694_ _6027_/CLK _5694_/D vssd1 vssd1 vccd1 vccd1 _5694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4645_ _5693_/Q _5670_/Q _4645_/S vssd1 vssd1 vccd1 vccd1 _4645_/X sky130_fd_sc_hd__mux2_1
X_4576_ _4575_/B _4574_/X _4575_/Y _4460_/X vssd1 vssd1 vccd1 vccd1 _5876_/D sky130_fd_sc_hd__o211a_1
X_3527_ _5864_/Q vssd1 vssd1 vccd1 vccd1 _3529_/A sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_39_wb_clk_i_A clkbuf_3_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3458_ _3158_/A _2863_/X _2885_/Y _3315_/Y _3457_/X vssd1 vssd1 vccd1 vccd1 _3489_/B
+ sky130_fd_sc_hd__a41o_1
X_3389_ _3389_/A _5281_/A _3066_/B vssd1 vssd1 vccd1 vccd1 _3407_/B sky130_fd_sc_hd__or3b_1
XFILLER_57_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5128_ _5145_/B vssd1 vssd1 vccd1 vccd1 _5138_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__4095__A _4095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5059_ _5059_/A vssd1 vssd1 vccd1 vccd1 _5059_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_72_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_36_wb_clk_i clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5929_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_48_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4430_ _5845_/Q _4429_/X _4433_/S vssd1 vssd1 vccd1 vccd1 _4431_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4731__A0 _6101_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3084__A _4466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6100_ _6138_/CLK _6100_/D vssd1 vssd1 vccd1 vccd1 _6100_/Q sky130_fd_sc_hd__dfxtp_1
X_4361_ _5824_/Q _4359_/X _4374_/S vssd1 vssd1 vccd1 vccd1 _4362_/A sky130_fd_sc_hd__mux2_1
X_4292_ _3354_/X _4322_/A _4243_/A vssd1 vssd1 vccd1 vccd1 _4294_/C sky130_fd_sc_hd__a21oi_1
X_3312_ _2950_/B _3312_/B _3312_/C _3312_/D vssd1 vssd1 vccd1 vccd1 _3326_/A sky130_fd_sc_hd__and4b_2
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6031_ _6031_/CLK _6031_/D vssd1 vssd1 vccd1 vccd1 _6031_/Q sky130_fd_sc_hd__dfxtp_1
X_3243_ _3243_/A _3243_/B _3243_/C _3243_/D vssd1 vssd1 vccd1 vccd1 _3244_/C sky130_fd_sc_hd__and4_1
XFILLER_66_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3174_ _5922_/Q vssd1 vssd1 vccd1 vccd1 _3174_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5815_ _6005_/CLK _5815_/D vssd1 vssd1 vccd1 vccd1 _5815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3259__A _3466_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2958_ _3429_/B _3424_/B vssd1 vssd1 vccd1 vccd1 _3476_/C sky130_fd_sc_hd__nor2_1
X_5746_ _6131_/CLK _5746_/D vssd1 vssd1 vccd1 vccd1 _5746_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3222__B1 _3221_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5677_ _5702_/CLK _5677_/D vssd1 vssd1 vccd1 vccd1 _5677_/Q sky130_fd_sc_hd__dfxtp_1
X_2889_ _3873_/C vssd1 vssd1 vccd1 vccd1 _3159_/B sky130_fd_sc_hd__clkbuf_2
X_4628_ _6115_/Q _4626_/X _4667_/S vssd1 vssd1 vccd1 vccd1 _4628_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4559_ _3139_/Y _5744_/Q _3509_/A vssd1 vssd1 vccd1 vccd1 _4559_/X sky130_fd_sc_hd__a21o_1
XFILLER_89_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4253__A2 _3826_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_470 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_378 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5384__A _5384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput61 _5888_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[75] sky130_fd_sc_hd__buf_2
Xoutput50 _5877_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[64] sky130_fd_sc_hd__buf_2
Xoutput72 _5899_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[86] sky130_fd_sc_hd__buf_2
XANTENNA__3632__A _3632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3930_ _3930_/A _3939_/A vssd1 vssd1 vccd1 vccd1 _3964_/A sky130_fd_sc_hd__nor2_1
XFILLER_63_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5278__B _5278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3861_ _3861_/A _3921_/B vssd1 vssd1 vccd1 vccd1 _3861_/X sky130_fd_sc_hd__and2_1
XFILLER_16_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3792_ _3966_/A _3792_/B vssd1 vssd1 vccd1 vccd1 _3793_/A sky130_fd_sc_hd__and2_1
X_5600_ _3582_/X _5580_/A _5599_/X _5597_/X vssd1 vssd1 vccd1 vccd1 _6104_/D sky130_fd_sc_hd__o211a_1
X_5531_ _6079_/Q _5533_/B vssd1 vssd1 vccd1 vccd1 _5531_/X sky130_fd_sc_hd__or2_1
XANTENNA__3807__A _4220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5462_ _5393_/X _5449_/X _5460_/X _5461_/X vssd1 vssd1 vccd1 vccd1 _6053_/D sky130_fd_sc_hd__o211a_1
X_5393_ _5393_/A vssd1 vssd1 vccd1 vccd1 _5393_/X sky130_fd_sc_hd__buf_2
X_4413_ _6063_/Q _5839_/Q _4426_/S vssd1 vssd1 vccd1 vccd1 _4413_/X sky130_fd_sc_hd__mux2_1
X_4344_ _5819_/Q _4341_/X _4357_/S vssd1 vssd1 vccd1 vccd1 _4345_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4275_ _5808_/Q _5807_/Q _4275_/C vssd1 vssd1 vccd1 vccd1 _4276_/C sky130_fd_sc_hd__and3_1
XFILLER_86_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4468__C1 _3331_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6014_ _6014_/CLK _6014_/D vssd1 vssd1 vccd1 vccd1 _6014_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3226_ _5933_/Q vssd1 vssd1 vccd1 vccd1 _3226_/Y sky130_fd_sc_hd__inv_2
X_3157_ _6123_/Q vssd1 vssd1 vccd1 vccd1 _4322_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_54_212 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3088_ _5256_/A vssd1 vssd1 vccd1 vccd1 _4237_/C sky130_fd_sc_hd__inv_2
XFILLER_54_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5729_ _5736_/CLK _5729_/D vssd1 vssd1 vccd1 vccd1 _5729_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5499__A1 _5353_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5379__A _5579_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5423__A1 _3614_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_51_wb_clk_i clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6024_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_5_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4458__A _4458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4060_ _4060_/A vssd1 vssd1 vccd1 vccd1 _5761_/D sky130_fd_sc_hd__clkbuf_1
X_3011_ _3836_/A vssd1 vssd1 vccd1 vccd1 _3375_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_91_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4962_ _4955_/X _4968_/C _4961_/X vssd1 vssd1 vccd1 vccd1 _4963_/B sky130_fd_sc_hd__a21bo_1
XFILLER_17_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3913_ _3913_/A _3913_/B _4473_/B vssd1 vssd1 vccd1 vccd1 _3914_/S sky130_fd_sc_hd__or3_1
X_4893_ _5967_/Q _4917_/B vssd1 vssd1 vccd1 vccd1 _4893_/X sky130_fd_sc_hd__or2_1
X_3844_ _5813_/Q _5228_/B _3844_/C _4438_/A vssd1 vssd1 vccd1 vccd1 _3845_/D sky130_fd_sc_hd__or4b_2
X_3775_ _3784_/A _3775_/B vssd1 vssd1 vccd1 vccd1 _3776_/A sky130_fd_sc_hd__and2_1
X_5514_ _5514_/A vssd1 vssd1 vccd1 vccd1 _5514_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5445_ _6048_/Q _5445_/B vssd1 vssd1 vccd1 vccd1 _5445_/X sky130_fd_sc_hd__or2_1
X_5376_ _5376_/A vssd1 vssd1 vccd1 vccd1 _5376_/X sky130_fd_sc_hd__buf_2
XANTENNA__5471__B _5471_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3272__A _4436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4327_ _4327_/A _4401_/B vssd1 vssd1 vccd1 vccd1 _4327_/Y sky130_fd_sc_hd__nor2_1
XFILLER_86_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4258_ _4256_/X _4257_/X _4259_/A vssd1 vssd1 vccd1 vccd1 _4258_/X sky130_fd_sc_hd__o21a_1
X_3209_ _5936_/Q vssd1 vssd1 vccd1 vccd1 _5012_/A sky130_fd_sc_hd__inv_2
XANTENNA__5653__A1 _5393_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4189_ _4189_/A vssd1 vssd1 vccd1 vccd1 _5798_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4916__A0 _5962_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3498__A3 _3497_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3560_ _5739_/Q vssd1 vssd1 vccd1 vccd1 _3561_/A sky130_fd_sc_hd__inv_2
X_5230_ _3874_/B _3872_/X _5229_/A vssd1 vssd1 vccd1 vccd1 _5230_/X sky130_fd_sc_hd__a21o_1
X_3491_ _4095_/A vssd1 vssd1 vccd1 vccd1 _3491_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4135__A1 _3037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5161_ _5062_/X _5149_/X _5160_/X _5158_/X vssd1 vssd1 vccd1 vccd1 _5982_/D sky130_fd_sc_hd__o211a_1
XFILLER_68_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4112_ _4112_/A vssd1 vssd1 vccd1 vccd1 _5776_/D sky130_fd_sc_hd__clkbuf_1
X_5092_ _5062_/X _5080_/X _5091_/X _5087_/X vssd1 vssd1 vccd1 vccd1 _5958_/D sky130_fd_sc_hd__o211a_1
XFILLER_83_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4043_ _4043_/A vssd1 vssd1 vccd1 vccd1 _5756_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3820__A _3820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5994_ _6002_/CLK _5994_/D vssd1 vssd1 vccd1 vccd1 _5994_/Q sky130_fd_sc_hd__dfxtp_1
X_4945_ _5981_/Q _4928_/B _4944_/Y _4940_/X vssd1 vssd1 vccd1 vccd1 _5917_/D sky130_fd_sc_hd__o211a_1
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4876_ _4870_/X _4873_/X _4874_/X _4875_/X vssd1 vssd1 vccd1 vccd1 _4876_/X sky130_fd_sc_hd__o211a_1
XFILLER_32_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3827_ _5241_/C _3901_/A _3826_/X vssd1 vssd1 vccd1 vccd1 _3828_/B sky130_fd_sc_hd__a21bo_1
X_3758_ _3758_/A vssd1 vssd1 vccd1 vccd1 _5702_/D sky130_fd_sc_hd__clkbuf_1
X_3689_ _3701_/A _3689_/B vssd1 vssd1 vccd1 vccd1 _3690_/A sky130_fd_sc_hd__and2_1
X_5428_ _5471_/B _5624_/B vssd1 vssd1 vccd1 vccd1 _5445_/B sky130_fd_sc_hd__nor2_1
XFILLER_87_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5359_ _5357_/X _5347_/X _5358_/X _5355_/X vssd1 vssd1 vccd1 vccd1 _6019_/D sky130_fd_sc_hd__o211a_1
XFILLER_59_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4062__A0 _6105_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xuser_proj_example_215 vssd1 vssd1 vccd1 vccd1 user_proj_example_215/HI la_data_out[122]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_237 vssd1 vssd1 vccd1 vccd1 user_proj_example_237/HI wbs_dat_o[16]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_226 vssd1 vssd1 vccd1 vccd1 user_proj_example_226/HI wbs_dat_o[5]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_204 vssd1 vssd1 vccd1 vccd1 user_proj_example_204/HI la_data_out[111]
+ sky130_fd_sc_hd__conb_1
XFILLER_11_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xuser_proj_example_259 vssd1 vssd1 vccd1 vccd1 io_out[7] user_proj_example_259/LO
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_248 vssd1 vssd1 vccd1 vccd1 user_proj_example_248/HI wbs_dat_o[27]
+ sky130_fd_sc_hd__conb_1
XFILLER_2_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5617__A1 _3611_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3628__A0 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2991_ _3435_/A _3350_/B _5304_/A vssd1 vssd1 vccd1 vccd1 _2991_/X sky130_fd_sc_hd__and3b_1
XFILLER_61_376 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4730_ _4781_/A vssd1 vssd1 vccd1 vccd1 _4771_/S sky130_fd_sc_hd__clkbuf_2
X_4661_ _6046_/Q _4654_/X _4610_/X _4660_/X vssd1 vssd1 vccd1 vccd1 _4661_/X sky130_fd_sc_hd__a211o_1
X_3612_ _5663_/Q _3618_/B vssd1 vssd1 vccd1 vccd1 _3612_/X sky130_fd_sc_hd__or2_1
X_4592_ _4883_/A vssd1 vssd1 vccd1 vccd1 _4781_/A sky130_fd_sc_hd__clkbuf_2
X_3543_ _4548_/A _5859_/Q _3540_/X _3556_/A _3408_/B vssd1 vssd1 vccd1 vccd1 _3544_/D
+ sky130_fd_sc_hd__a311o_1
XANTENNA_clkbuf_leaf_29_wb_clk_i_A clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3474_ _3482_/A _3869_/A _3870_/A _3829_/D _3287_/X vssd1 vssd1 vccd1 vccd1 _3474_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_88_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5213_ _5062_/A _6000_/Q _5216_/S vssd1 vssd1 vccd1 vccd1 _5214_/B sky130_fd_sc_hd__mux2_1
X_5144_ _5072_/X _5125_/A _5143_/X _5141_/X vssd1 vssd1 vccd1 vccd1 _5977_/D sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_0_wb_clk_i_A wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5075_ _5075_/A vssd1 vssd1 vccd1 vccd1 _5075_/X sky130_fd_sc_hd__clkbuf_2
X_4026_ _4026_/A vssd1 vssd1 vccd1 vccd1 _5751_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5977_ _5986_/CLK _5977_/D vssd1 vssd1 vccd1 vccd1 _5977_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5477__A _5529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4928_ _4928_/A _4928_/B vssd1 vssd1 vccd1 vccd1 _4928_/Y sky130_fd_sc_hd__nand2_1
XFILLER_60_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4859_ _4859_/A vssd1 vssd1 vccd1 vccd1 _4859_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_502 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5387__A _5387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3190_ _5923_/Q _5914_/Q vssd1 vssd1 vccd1 vccd1 _3190_/X sky130_fd_sc_hd__or2_1
XFILLER_78_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4466__A _4466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5900_ _6088_/CLK _5900_/D vssd1 vssd1 vccd1 vccd1 _5900_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5831_ _6050_/CLK _5831_/D vssd1 vssd1 vccd1 vccd1 _5831_/Q sky130_fd_sc_hd__dfxtp_1
X_2974_ _2997_/A vssd1 vssd1 vccd1 vccd1 _3826_/C sky130_fd_sc_hd__buf_2
X_5762_ _6018_/CLK _5762_/D vssd1 vssd1 vccd1 vccd1 _5762_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4713_ _6051_/Q _4706_/X _4664_/X _4712_/X vssd1 vssd1 vccd1 vccd1 _4713_/X sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_6_wb_clk_i clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6067_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_5693_ _6067_/CLK _5693_/D vssd1 vssd1 vccd1 vccd1 _5693_/Q sky130_fd_sc_hd__dfxtp_1
X_4644_ _5880_/Q _4579_/X _4642_/X _4643_/X vssd1 vssd1 vccd1 vccd1 _5880_/D sky130_fd_sc_hd__a22o_1
X_4575_ _4575_/A _4575_/B vssd1 vssd1 vccd1 vccd1 _4575_/Y sky130_fd_sc_hd__nand2_1
X_3526_ _4450_/B _4331_/B _3412_/X _3935_/C vssd1 vssd1 vccd1 vccd1 _6127_/D sky130_fd_sc_hd__a22o_1
XFILLER_89_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3457_ _3454_/X _3304_/B _3326_/A _3455_/X _3456_/X vssd1 vssd1 vccd1 vccd1 _3457_/X
+ sky130_fd_sc_hd__a41o_1
X_3388_ _6125_/Q vssd1 vssd1 vccd1 vccd1 _5249_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5127_ _5471_/B _5150_/B vssd1 vssd1 vccd1 vccd1 _5145_/B sky130_fd_sc_hd__nor2_1
XFILLER_57_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5058_ _5056_/X _5050_/X _5057_/X _5043_/X vssd1 vssd1 vccd1 vccd1 _5948_/D sky130_fd_sc_hd__o211a_1
XFILLER_84_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4009_ _5284_/A _3925_/Y _3522_/B vssd1 vssd1 vccd1 vccd1 _5747_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__5462__C1 _5461_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3439__B _5327_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4050__S _4063_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input32_A la_data_in[57] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3349__B _3854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4360_ _4397_/S vssd1 vssd1 vccd1 vccd1 _4374_/S sky130_fd_sc_hd__clkbuf_2
X_3311_ _4438_/B vssd1 vssd1 vccd1 vccd1 _3483_/B sky130_fd_sc_hd__clkbuf_2
X_4291_ _3842_/B _4291_/B _4291_/C _4291_/D vssd1 vssd1 vccd1 vccd1 _4297_/B sky130_fd_sc_hd__and4b_2
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6030_ _6031_/CLK _6030_/D vssd1 vssd1 vccd1 vccd1 _6030_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3242_ _5387_/A _5928_/Q _4986_/B _5384_/A _3241_/X vssd1 vssd1 vccd1 vccd1 _3243_/D
+ sky130_fd_sc_hd__a221oi_1
X_3173_ _5915_/Q vssd1 vssd1 vccd1 vccd1 _4939_/A sky130_fd_sc_hd__inv_2
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3470__A1 _3469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5814_ _6005_/CLK _5814_/D vssd1 vssd1 vccd1 vccd1 _5814_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2957_ _3400_/B vssd1 vssd1 vccd1 vccd1 _3424_/B sky130_fd_sc_hd__clkbuf_2
X_5745_ _6121_/CLK hold1/X vssd1 vssd1 vccd1 vccd1 _5745_/Q sky130_fd_sc_hd__dfxtp_1
X_2888_ _5812_/Q _5811_/Q _5810_/Q _5809_/Q vssd1 vssd1 vccd1 vccd1 _3873_/C sky130_fd_sc_hd__or4bb_2
X_5676_ _5702_/CLK _5676_/D vssd1 vssd1 vccd1 vccd1 _5676_/Q sky130_fd_sc_hd__dfxtp_1
X_4627_ _4779_/A vssd1 vssd1 vccd1 vccd1 _4667_/S sky130_fd_sc_hd__clkbuf_2
X_4558_ _4558_/A vssd1 vssd1 vccd1 vccd1 _5871_/D sky130_fd_sc_hd__clkbuf_1
X_4489_ _5847_/Q _4489_/B vssd1 vssd1 vccd1 vccd1 _4489_/Y sky130_fd_sc_hd__nand2_1
X_3509_ _3509_/A _3509_/B _3954_/A vssd1 vssd1 vccd1 vccd1 _3509_/X sky130_fd_sc_hd__and3_1
XFILLER_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3213__A1 _6023_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3213__B2 _6017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3884__S _4041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput51 _5878_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[65] sky130_fd_sc_hd__buf_2
Xoutput62 _5889_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[76] sky130_fd_sc_hd__buf_2
Xoutput73 _5900_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[87] sky130_fd_sc_hd__buf_2
XANTENNA__3819__A3 _4331_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4744__A _5403_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3860_ _3874_/B _3897_/D vssd1 vssd1 vccd1 vccd1 _3921_/B sky130_fd_sc_hd__or2_1
X_3791_ _3617_/A _5712_/Q _3791_/S vssd1 vssd1 vccd1 vccd1 _3792_/B sky130_fd_sc_hd__mux2_1
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5530_ _5396_/X _5514_/A _5528_/X _5529_/X vssd1 vssd1 vccd1 vccd1 _6078_/D sky130_fd_sc_hd__o211a_1
XANTENNA__3807__B _3928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5461_ _5461_/A vssd1 vssd1 vccd1 vccd1 _5461_/X sky130_fd_sc_hd__buf_2
X_4412_ _4432_/S vssd1 vssd1 vccd1 vccd1 _4426_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__4704__A1 _5886_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5392_ _5389_/X _5378_/X _5390_/X _5391_/X vssd1 vssd1 vccd1 vccd1 _6028_/D sky130_fd_sc_hd__o211a_1
X_4343_ _4397_/S vssd1 vssd1 vccd1 vccd1 _4357_/S sky130_fd_sc_hd__clkbuf_2
X_4274_ _5807_/Q _4275_/C _5808_/Q vssd1 vssd1 vccd1 vccd1 _4276_/B sky130_fd_sc_hd__a21oi_1
XFILLER_59_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3225_ _5855_/Q vssd1 vssd1 vccd1 vccd1 _4982_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6013_ _6014_/CLK _6013_/D vssd1 vssd1 vccd1 vccd1 _6013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3156_ _5544_/A vssd1 vssd1 vccd1 vccd1 _3632_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_27_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3087_ _6132_/Q vssd1 vssd1 vccd1 vccd1 _5256_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_54_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4654__A _4706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5469__B _5469_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3989_ _3989_/A vssd1 vssd1 vccd1 vccd1 _5733_/D sky130_fd_sc_hd__clkbuf_1
X_5728_ _5808_/CLK _5728_/D vssd1 vssd1 vccd1 vccd1 _5728_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4943__A1 _5980_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5659_ _6108_/CLK _5659_/D vssd1 vssd1 vccd1 vccd1 _5659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5379__B _5379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4934__A1 _6038_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_20_wb_clk_i _5836_/CLK vssd1 vssd1 vccd1 vccd1 _6131_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_output63_A _5890_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3010_ _3469_/B _3010_/B _3017_/B vssd1 vssd1 vccd1 vccd1 _3022_/C sky130_fd_sc_hd__and3_1
XFILLER_76_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4961_ _5920_/Q _4958_/B _5921_/Q vssd1 vssd1 vccd1 vccd1 _4961_/X sky130_fd_sc_hd__a21o_1
XFILLER_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3912_ _5234_/B _3886_/B _3921_/C _3861_/X vssd1 vssd1 vccd1 vccd1 _4473_/B sky130_fd_sc_hd__o211ai_2
X_4892_ _5959_/Q _4891_/X _4916_/S vssd1 vssd1 vccd1 vccd1 _4892_/X sky130_fd_sc_hd__mux2_1
X_3843_ _4002_/A _3843_/B vssd1 vssd1 vccd1 vccd1 _4283_/C sky130_fd_sc_hd__nand2_1
XFILLER_32_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3774_ _3601_/A _5707_/Q _3780_/S vssd1 vssd1 vccd1 vccd1 _3775_/B sky130_fd_sc_hd__mux2_1
X_5513_ _5579_/A _5535_/B vssd1 vssd1 vccd1 vccd1 _5514_/A sky130_fd_sc_hd__or2_1
X_5444_ _5369_/X _5427_/A _5443_/X _5435_/X vssd1 vssd1 vccd1 vccd1 _6047_/D sky130_fd_sc_hd__o211a_1
XANTENNA__3553__A _3553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5375_ _5373_/X _5354_/B _5374_/X _5371_/X vssd1 vssd1 vccd1 vccd1 _6024_/D sky130_fd_sc_hd__o211a_1
XANTENNA__3272__B _3272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4326_ _3494_/A _3484_/B _3800_/Y vssd1 vssd1 vccd1 vccd1 _4401_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__3900__A2 _3821_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4257_ _3858_/A _3264_/A _3042_/X vssd1 vssd1 vccd1 vccd1 _4257_/X sky130_fd_sc_hd__o21a_1
XFILLER_86_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3208_ _5937_/Q vssd1 vssd1 vccd1 vccd1 _3208_/Y sky130_fd_sc_hd__inv_2
X_4188_ _5798_/Q _4186_/X _4200_/S vssd1 vssd1 vccd1 vccd1 _4189_/A sky130_fd_sc_hd__mux2_1
X_3139_ _4529_/A vssd1 vssd1 vccd1 vccd1 _3139_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_514 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3416__A1 _3272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_128 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3129__B_N _5713_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3463__A _3481_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_19_wb_clk_i_A _5836_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3490_ _4113_/A vssd1 vssd1 vccd1 vccd1 _4095_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__5332__A1 _6065_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3894__A1 _3880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5160_ _5982_/Q _5162_/B vssd1 vssd1 vccd1 vccd1 _5160_/X sky130_fd_sc_hd__or2_1
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3894__B2 _5768_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4111_ _5776_/Q _4110_/X _4116_/S vssd1 vssd1 vccd1 vccd1 _4112_/A sky130_fd_sc_hd__mux2_1
X_5091_ _5958_/Q _5093_/B vssd1 vssd1 vccd1 vccd1 _5091_/X sky130_fd_sc_hd__or2_1
X_4042_ _5756_/Q _4041_/X _4046_/S vssd1 vssd1 vccd1 vccd1 _4043_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5993_ _6002_/CLK _5993_/D vssd1 vssd1 vccd1 vccd1 _5993_/Q sky130_fd_sc_hd__dfxtp_1
X_4944_ _4944_/A _4944_/B vssd1 vssd1 vccd1 vccd1 _4944_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_58_wb_clk_i_A clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4875_ _5126_/A vssd1 vssd1 vccd1 vccd1 _4875_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3826_ _4281_/A _4217_/A _3826_/C vssd1 vssd1 vccd1 vccd1 _3826_/X sky130_fd_sc_hd__or3_1
XANTENNA__3267__B _3928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3757_ _3768_/A _3757_/B vssd1 vssd1 vccd1 vccd1 _3758_/A sky130_fd_sc_hd__and2_1
X_3688_ _3598_/A _5683_/Q _3697_/S vssd1 vssd1 vccd1 vccd1 _3689_/B sky130_fd_sc_hd__mux2_1
X_5427_ _5427_/A vssd1 vssd1 vccd1 vccd1 _5427_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5358_ _6019_/Q _5367_/B vssd1 vssd1 vccd1 vccd1 _5358_/X sky130_fd_sc_hd__or2_1
X_4309_ _5811_/Q _4309_/B vssd1 vssd1 vccd1 vccd1 _4309_/X sky130_fd_sc_hd__xor2_1
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5289_ _5289_/A _5289_/B vssd1 vssd1 vccd1 vccd1 _5289_/Y sky130_fd_sc_hd__nor2_1
XFILLER_74_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4842__A _4842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4062__A1 _3869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4053__S _4063_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_proj_example_216 vssd1 vssd1 vccd1 vccd1 user_proj_example_216/HI la_data_out[123]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_227 vssd1 vssd1 vccd1 vccd1 user_proj_example_227/HI wbs_dat_o[6]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_205 vssd1 vssd1 vccd1 vccd1 user_proj_example_205/HI la_data_out[112]
+ sky130_fd_sc_hd__conb_1
XFILLER_23_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuser_proj_example_249 vssd1 vssd1 vccd1 vccd1 user_proj_example_249/HI wbs_dat_o[28]
+ sky130_fd_sc_hd__conb_1
Xuser_proj_example_238 vssd1 vssd1 vccd1 vccd1 user_proj_example_238/HI wbs_dat_o[17]
+ sky130_fd_sc_hd__conb_1
XFILLER_78_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3628__A1 _5666_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2990_ _5277_/C _2990_/B vssd1 vssd1 vccd1 vccd1 _5304_/A sky130_fd_sc_hd__nor2_1
XFILLER_64_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3368__A _3897_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4660_ _4611_/X _4658_/X _4659_/X _4620_/X vssd1 vssd1 vccd1 vccd1 _4660_/X sky130_fd_sc_hd__o211a_1
X_3611_ _3611_/A vssd1 vssd1 vccd1 vccd1 _3611_/X sky130_fd_sc_hd__clkbuf_2
X_4591_ _4594_/A _4591_/B _4594_/C vssd1 vssd1 vccd1 vccd1 _4883_/A sky130_fd_sc_hd__or3_2
XANTENNA__5583__A _6097_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3542_ _3542_/A vssd1 vssd1 vccd1 vccd1 _3556_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3473_ _5241_/C vssd1 vssd1 vccd1 vccd1 _3869_/A sky130_fd_sc_hd__clkbuf_2
X_5212_ _5212_/A vssd1 vssd1 vccd1 vccd1 _5999_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5143_ _5977_/Q _5145_/B vssd1 vssd1 vccd1 vccd1 _5143_/X sky130_fd_sc_hd__or2_1
XANTENNA__3831__A _5250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5074_ _5072_/X _5050_/A _5073_/X _5067_/X vssd1 vssd1 vccd1 vccd1 _5953_/D sky130_fd_sc_hd__o211a_1
X_4025_ _5751_/Q _4024_/X _4028_/S vssd1 vssd1 vccd1 vccd1 _4026_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5976_ _5986_/CLK _5976_/D vssd1 vssd1 vccd1 vccd1 _5976_/Q sky130_fd_sc_hd__dfxtp_1
X_4927_ _4927_/A vssd1 vssd1 vccd1 vccd1 _4928_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4858_ _4858_/A vssd1 vssd1 vccd1 vccd1 _4858_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3809_ _3405_/A _3497_/X _3849_/C _3405_/X _5835_/Q vssd1 vssd1 vccd1 vccd1 _3809_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_20_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4789_ _5660_/Q _4788_/X _4821_/S vssd1 vssd1 vccd1 vccd1 _4789_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3741__A _3750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_406 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4572__A _5186_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_160 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5830_ _6050_/CLK _5830_/D vssd1 vssd1 vccd1 vccd1 _5830_/Q sky130_fd_sc_hd__dfxtp_1
X_2973_ _3440_/A _3820_/B _3360_/B _2972_/X vssd1 vssd1 vccd1 vccd1 _2973_/X sky130_fd_sc_hd__a31o_1
XFILLER_61_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5761_ _6005_/CLK _5761_/D vssd1 vssd1 vccd1 vccd1 _5761_/Q sky130_fd_sc_hd__dfxtp_1
X_4712_ _4665_/X _4710_/X _4711_/X _4670_/X vssd1 vssd1 vccd1 vccd1 _4712_/X sky130_fd_sc_hd__o211a_1
X_5692_ _5941_/CLK _5692_/D vssd1 vssd1 vccd1 vccd1 _5692_/Q sky130_fd_sc_hd__dfxtp_1
X_4643_ _6020_/Q _4606_/X _4607_/X vssd1 vssd1 vccd1 vccd1 _4643_/X sky130_fd_sc_hd__o21a_1
X_4574_ _4567_/Y _3147_/B _4529_/A vssd1 vssd1 vccd1 vccd1 _4574_/X sky130_fd_sc_hd__o21a_1
X_3525_ _3525_/A vssd1 vssd1 vccd1 vccd1 _4331_/B sky130_fd_sc_hd__clkbuf_2
X_3456_ _2899_/A _3047_/X _3042_/X _3037_/Y _3412_/A vssd1 vssd1 vccd1 vccd1 _3456_/X
+ sky130_fd_sc_hd__a41o_1
X_3387_ _3387_/A vssd1 vssd1 vccd1 vccd1 _6121_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5126_ _5126_/A vssd1 vssd1 vccd1 vccd1 _5471_/B sky130_fd_sc_hd__buf_2
XFILLER_29_127 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5057_ _5948_/Q _5066_/B vssd1 vssd1 vccd1 vccd1 _5057_/X sky130_fd_sc_hd__or2_1
X_4008_ _4008_/A vssd1 vssd1 vccd1 vccd1 _5746_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5488__A _5529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5959_ _5959_/CLK _5959_/D vssd1 vssd1 vccd1 vccd1 _5959_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3736__A _3750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input25_A la_data_in[50] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_45_wb_clk_i clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5986_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_45_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5508__A1 _5366_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3310_ _3462_/C _3310_/B vssd1 vssd1 vccd1 vccd1 _3310_/X sky130_fd_sc_hd__or2_1
X_4290_ _3802_/B _3367_/Y _3830_/B _4288_/Y _4289_/Y vssd1 vssd1 vccd1 vccd1 _4291_/D
+ sky130_fd_sc_hd__o2111a_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3241_ _6028_/Q _5929_/Q vssd1 vssd1 vccd1 vccd1 _3241_/X sky130_fd_sc_hd__xor2_1
X_3172_ _5853_/Q vssd1 vssd1 vccd1 vccd1 _4946_/C sky130_fd_sc_hd__clkbuf_2
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5813_ _5813_/CLK _5813_/D vssd1 vssd1 vccd1 vccd1 _5813_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2956_ _2928_/Y _5289_/A _2948_/X _2955_/X vssd1 vssd1 vccd1 vccd1 _3022_/A sky130_fd_sc_hd__o31a_1
X_5744_ _6121_/CLK _5744_/D vssd1 vssd1 vccd1 vccd1 _5744_/Q sky130_fd_sc_hd__dfxtp_1
X_2887_ _3839_/B vssd1 vssd1 vccd1 vccd1 _3480_/B sky130_fd_sc_hd__buf_2
X_5675_ _6080_/CLK _5675_/D vssd1 vssd1 vccd1 vccd1 _5675_/Q sky130_fd_sc_hd__dfxtp_1
X_4626_ _5691_/Q _5668_/Q _4645_/S vssd1 vssd1 vccd1 vccd1 _4626_/X sky130_fd_sc_hd__mux2_1
X_4557_ _3454_/X _4554_/X _4557_/S vssd1 vssd1 vccd1 vccd1 _4558_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4488_ _4488_/A vssd1 vssd1 vccd1 vccd1 _4489_/B sky130_fd_sc_hd__inv_2
X_3508_ _3929_/B _3508_/B _3508_/C vssd1 vssd1 vccd1 vccd1 _3954_/A sky130_fd_sc_hd__and3_1
XFILLER_77_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3439_ _3439_/A _5327_/B _3870_/A vssd1 vssd1 vccd1 vccd1 _3440_/D sky130_fd_sc_hd__and3_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5109_ _5964_/Q _5116_/B vssd1 vssd1 vccd1 vccd1 _5109_/X sky130_fd_sc_hd__or2_1
XFILLER_57_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6089_ _6115_/CLK _6089_/D vssd1 vssd1 vccd1 vccd1 _6089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput52 _5879_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[66] sky130_fd_sc_hd__buf_2
Xoutput74 _5901_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[88] sky130_fd_sc_hd__buf_2
Xoutput63 _5890_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[77] sky130_fd_sc_hd__buf_2
XFILLER_0_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3790_ _3790_/A vssd1 vssd1 vccd1 vccd1 _5711_/D sky130_fd_sc_hd__clkbuf_1
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5460_ _6053_/Q _5460_/B vssd1 vssd1 vccd1 vccd1 _5460_/X sky130_fd_sc_hd__or2_1
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4411_ _4411_/A vssd1 vssd1 vccd1 vccd1 _5839_/D sky130_fd_sc_hd__clkbuf_1
X_5391_ _5391_/A vssd1 vssd1 vccd1 vccd1 _5391_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4342_ _4366_/A _3406_/Y _3812_/S vssd1 vssd1 vccd1 vccd1 _4397_/S sky130_fd_sc_hd__a21oi_4
X_4273_ _4273_/A vssd1 vssd1 vccd1 vccd1 _5807_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4580__B_N _3564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6012_ _6012_/CLK _6012_/D vssd1 vssd1 vccd1 vccd1 _6012_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4000__A _5188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3224_ _3218_/X _3215_/C _5012_/B vssd1 vssd1 vccd1 vccd1 _3224_/Y sky130_fd_sc_hd__a21oi_1
.ends

